af
arkeo
astro
av
be
bi
bio
cyklo
e
elektro
engångs
er
ex
femto
fort
frilufts
fysio
för
geo
gyneko
gôr
huvud
justitie
kata
kontra
kosmo
lexiko
medel
mid
mikro
o
paleo
pseudo
psyko
re
riks
sam
styv
svär
sär
tele
toxiko
tri
van
veder
ärke
örlogs
över
