a
aktig
al
an
ande
ar
are
arie
arna
ast
atör
bar
bo
d
dd
de
dimensionell
dom
e
ell
else
en
ende
er
era
eri
erna
erska
es
et
faldig
falt
gnos
graf
grafi
gram
het
huvud
i
ier
ifiera
ig
ing
inna
is
isera
isk
it
itet
iv
ledes
lig
log
logi
lunda
lös
makare
mang
ment
mässig
n
na
ne
ning
nomi
or
orna
r
re
rna
s
sam
sel
sk
skap
son
städes
t
te
tion
ur
vis
är
ör
ös
