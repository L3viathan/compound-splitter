      4 []
      1 [���]
      2 ]
    518 �
     26 ��
     23 ���
      8 ����
      2 �����
      1 ������
      3 �������
      1 ��������
      3 ����������
      3 �����������
      1 ������������
    208 a
      1 [a�]
     33 å
     13 Å
      1 ä
      2 Ä
      4 aa
      2 aaa
      4 aad
      2 aaföreningar
      1 aagenaes
      1 aagen�s
      1 aagrupper
      1 aai
      1 aal
      1 aantigenen
      1 aarhus
      3 aaron
     30 ab
      1 abaptiston
      1 abasi
      1 abbasid
      1 abbaye
      1 abbe
      1 abbey
      1 abborrverket
      1 abchazien
      1 abdominell
      4 abdominis
      1 abductionfenomenet
      1 abelius
      1 åberopas
      2 abilify
      1 ability
      1 abiogenes
      1 abiogenesiska
      3 ablation
      1 ablationsbehandling
      2 ablefari
      5 abnorm
      5 abnorma
      1 abnormala
      1 abnormalitet
      7 abnormaliteter
      3 abnormalt
      7 abnormt
      1 abo
      1 Åbo
      1 Åbolands
      1 aboriginer
      1 aboriginspråk
      1 abormaliteter
     73 abort
      1 abortansökan
      1 abortdagen
      9 aborten
     36 aborter
      1 aborteras
      2 abortering
      1 abortfrågan
      1 abortframkallande
      2 abortingrepp
      2 abortion
      1 abortivägg
      1 abortkritiker
      1 abortlag
      1 abortlagen
      1 abortlagstiftning
      1 abortmedel
      1 abortmetod
      1 abortmetoder
      1 abortmöjlighet
      2 abortpiller
      1 abortrådgivning
      1 abosystemet
      2 about
      1 aboutalib
      1 above
      2 abpa
      2 abraham
      1 abrahamitiska
      2 abram
      5 abrupt
      1 abrupta
      1 abs
      1 abscensanfall
      5 abscess
      2 abscessbildning
      3 abscessen
     13 abscesser
      2 absence
      1 absenor
      3 absens
      1 absensanfall
      2 absenser
      2 absentia
      1 abs�ns
     24 absolut
      9 absoluta
      1 absolutely
      1 absoluteras
      1 absolutionen
     13 absorbera
      5 absorberad
      2 absorberade
      1 absorberades
      5 absorberande
      8 absorberar
     18 absorberas
      2 absorberats
      1 absorbering
      4 absorption
      4 absorptionen
      1 absorptionsförmåga
      1 absorptionsgrad
      2 absorptionsyta
      2 absorptionsytan
      1 absorptiva
     10 abstinens
      2 abstinensbehandling
      5 abstinensbesvär
      1 abstinensen
      1 abstinensepilepsi
      1 abstinensepileptiska
      1 abstinensfas
      1 abstinensfenomen
      2 abstinenskomplikationer
      4 abstinenskramper
      1 abstinensliknande
      1 abstinent
      9 abstrakt
      2 abstrakta
      1 abstraktioner
      2 absurda
      1 absurdum
      7 absystemet
      1 absystemets
      2 abtoxin
      1 abtoxiner
      2 abtoxinet
      1 abu
      1 abvr
      2 ac
      2 aca
      2 acacia
      1 academic
      2 académie
      4 academy
      1 acanthamoeba
      2 acanthosis
      1 accelerationsnod
      1 accelerationsröret
      1 accelerationsspänningen
      1 accelerato
      1 accelerera
      1 accelererad
      2 accelererar
      6 accelereras
      1 accenten
      1 accentuation
      1 accentuerade
      2 accentueras
      1 accentueringsförsök
      6 acceptabel
      5 acceptabelt
      2 acceptabla
      4 acceptance
      4 acceptans
      3 acceptansen
      1 acceptens
      9 acceptera
      8 accepterad
      8 accepterade
      2 accepterades
      2 accepterar
      2 accepteras
     11 accepterat
      1 accepterats
      1 accepts
      1 accesorisk
      1 accessible
      1 accessoarer
      2 accessoriska
      1 accessorius
      1 according
      3 accumbenskärnan
      1 accumbensområdet
      1 accuminata
      4 ace
      2 acedia
      1 acefat
      1 aceh
      4 acehämmare
      1 acehämmarna
      2 acen
      2 acerebri
      1 aceruloplasminemi
      6 acetaldehyd
      1 acet�aldehyd�dehydrogenas
      1 acetaminofenparacetamol
      2 acetaminophen
      1 acetat
      1 acetatbågarna
      1 acetazolamid
      8 aceton
      1 acetonfria
      1 acetonliknande
      1 acetontricykloperoxid
      1 acetyl
      2 acetylcoa
      1 acetylcoakarboxylas
      1 acetylen
     16 acetylkolin
      2 acetylkolinesteras
      1 acetylkolinet
      1 acetylkolinreceptorer
      1 acetylkolinreceptorn
      1 acetylsalicylic
     14 acetylsalicylsyra
      1 acetylsalicylsyrapreparat
      1 achim
      7 acid
      1 acidofilusbakterier
      1 acidophilus
     25 acidos
      1 acidosen
      1 acids
      3 aciklovir
      1 acinosa
      1 äckla
      5 acklimatisering
      3 ackommodation
      1 ackommodationen
      1 ackommodationsförmågan
      1 ackommodationskraften
      2 ackommodationsvila
      2 ackommodera
      3 ackompanjemang
      1 ackoppling
      1 ackrediterade
      1 ackumulatorer
      1 ackumulera
      1 ackumulerar
      3 ackumuleras
      2 ackumulering
      2 ackumuleringen
      1 ackuschörska
      2 acne
      1 acokanthera
      3 aconitum
      1 acquired
      3 acrbr
      1 acre
      1 acrosin
      4 act
      1 acta
      1 actaea
      5 acth
      1 acthadenom
      1 actilyse
      1 actinobacillus
      1 actinomycetales
      1 actionhjältinna
      1 activated
      1 active
      1 activity
      2 acupuncture
      1 acus
      1 acuta
      4 acute
      1 acutifolius
      1 acwpolysackaridvacciner
      1 acwy
      1 acylgrupp
      4 ad
      2 ada
      1 Ådalen
      1 adam
      1 adamantan
      5 adams
      2 adamsstokes
      3 adaptation
      1 adapter
      3 adaption
      2 adaptiv
      9 adaptiva
      3 adaptivt
      6 add
      1 adderas
      1 addis
      2 addisons
      1 addisonschilder
      1 additativt
      1 addressed
      1 addressing
      2 adductus
      1 addukterna
      2 ade
     17 adekvat
      4 adekvata
      1 adel
      2 adelen
      1 ädelgasen
      1 adelmann
      1 ädelmetall
      1 ädelmetaller
      1 ädelröta
      1 Ädelröta
      1 ädelrötade
      2 adelsman
      1 adelsmän
      1 adelsmännen
      2 ädelsöta
      1 adelsrytteriets
      2 ädelsten
      1 ädelstenar
      2 adenin
      1 adenit
     12 adenocarcinom
      1 adenocarcinomtyp
      6 adenohypofysen
      1 adenoid
      1 adenoida
     12 adenom
      1 adenomet
      1 adenomvariant
      1 adenomyos
      2 adenosarkom
     10 adenosin
      1 adenosindeaminastest
      1 adenosindifosfat
      1 adenosindifosfatet
      1 adenosinreceptorer
      2 adenosintrifosfat
      5 adenovirus
      1 adenylatcyklas
     15 åderbråck
      3 Åderbråck
      1 åderbråckskirurgi
      1 åderbråcksvener
      2 åderförfettning
      1 Åderförfettning
      9 åderförkalkning
      1 åderförkalkningen
      1 åderförkalkningsplacken
      2 åderhinnan
      1 åderkalkade
      1 åderlåtas
     17 åderlåtning
      2 Åderlåtning
      1 Åderlåtningsmannen
      7 adh
      1 adhcc
     85 adhd
      6 adhdc
      1 adhdcoacher
      1 adhdcproblematik
      1 adhdfall
      2 adhdh
      1 adhdhjärnstruktur
      9 adhdi
      1 adhdigruppen
      1 adhdigrupperna
      1 adhdkombinerad
      1 adhdliknande
      1 adhdpi
      1 adhdproblematik
      1 adhdsymtom
      1 adhdvarianterna
      1 adherence
      1 adherencer
      1 adherens
      8 adherenser
      1 adhesiner
      2 adhesion
      1 adhesioner
      1 adhhalterna
      1 adhsekretion
      1 adipinsyra
      3 adipocyter
      1 adipocytokiner
      1 adipocytokinerna
      1 adiponektin
      1 adiposis
      2 adir
      1 adjektiv
      1 adjektivet
      3 adjuvans
      2 adjuvant
      2 adjuvantbehandling
      1 adl
      1 ädla
      1 ädle
      1 adliga
      1 administering
      1 administratiion
     11 administration
      1 administrationstid
      1 administrativ
      3 administrativa
      2 administrativt
      3 administrera
      1 administrerades
     11 administreras
      2 administrerats
      2 administrering
      1 administreringsform
      2 adolescens
      6 adolescensen
      3 adolescensens
      1 adolescere
      1 adolesent
      9 adolf
      1 adom
      1 adomvandlare
      2 adonis
      2 adonisarter
      1 adoptera
      1 adopterades
      1 adoption
      2 ados
      1 adr
      4 ådragit
      1 adramytes
      2 ådrar
      1 ådras
      1 adrenal
     39 adrenalin
      1 adrenalinliknande
      1 adrenalinutsöndring
      2 adrenerga
      2 adrenogenitalt
      2 adrenokortikotropiskt
      2 adrenokortikotropt
      1 adrenoleukodystrofi
      1 adrenomedullin
      1 adrenomyeloneuropati
      1 adressera
      1 adresserandet
      1 adrian
      1 ådrig
      3 ådror
      1 ådrorna
      1 ådrornas
      2 adsorberas
      8 adult
      3 adulta
      1 adults
      1 advaita
      2 advance
      1 advanced
      1 adventivrot
      1 adventivrotsbildning
      3 adventivrötter
      1 adventure
      2 adverse
      1 advokat
      1 advokater
      1 ae
      1 a�e
      1 aebelholt
     11 aedes
      1 aedesmyggor
      5 aegypti
      1 aemula
      1 aequalia
      1 aequalibus
      8 aerob
      5 aeroba
      1 aerobicspass
      1 aerobiska
      1 aerobt
      4 aerosol
      3 aerosoler
      1 aerosolsmitta
      1 aerosystems
      1 aerotolerant
      1 aeruginosa
      5 aesculapius
      1 aestivalis
      1 aeternitas
      1 aetheroleum
      1 aethiopica
      1 aethusa
      1 aex
      6 af
      1 afaki
     38 afasi
      1 afasidiagnoserna
      2 afasidrabbade
      1 afasier
      1 afasin
      1 afasisymptomen
      1 afasisymtom
      1 afasisyndrom
      1 afasityp
      1 affär
      2 affären
      3 affärer
      1 affärerna
      1 affärslivet
      2 affärsmän
      1 affärsområden
      1 affärsplan
      2 affärsverksamhet
      9 affekt
      2 affekter
      2 affekterna
      1 affektinkontinens
     12 affektiv
     21 affektiva
      1 affektivaperceptuella
      3 affektivt
      1 affiliering
      1 affinis
     15 affinitet
      2 affiniteten
      1 affinitetsmognad
      2 afghanistan
      1 afil
      1 afilter
      1 afiltret
      1 aflägsna
      4 afoni
      1 afoniröstavbrott
      1 afp
      1 africanum
     92 afrika
      1 afrikaner
      2 afrikansk
      7 afrikanska
      2 afrikanskt
      4 afrikas
      1 afroamerikaner
      2 afrodisiakum
      4 afs
      1 afsset
     10 afte
      1 aftershave
      1 aftonen
      1 aftonklänning
      1 aftonklänningar
      1 aftös
      1 aftösa
      1 äfwen
      1 afylaxi
      1 afzelii
      1 ag
      5 aga
      7 äga
      2 against
      1 agalactiae
      1 agamer
      5 ägare
      2 Ägare
      3 ägaren
      2 ägarens
      1 agaricaceae
      1 agaricus
      1 ägarnas
      1 ägas
      6 agave
      1 agavearter
      1 agavesläktet
      1 agavesläktets
      1 ägcellens
      2 ägda
     10 ägde
      1 age
      2 agence
      4 agency
      1 agendor
      2 agenesi
      3 agens
      2 agenset
      3 agent
      4 agenter
      1 agentur
      1 agenturer
     19 äger
     11 agera
      3 agerade
      3 agerande
      1 ageranden
     11 agerar
      1 ageratina
      2 ageratum
      1 agere
      1 agerörelsen
      3 ageusi
    124 ägg
      1 Ägg
      1 ägganlag
      1 ägganlagen
      2 äggblåsa
      1 äggblåsan
      1 äggblåsor
      1 äggblåsorna
     10 äggcell
     13 äggcellen
      2 Äggcellen
      3 äggcellens
     13 äggceller
      5 äggcellerna
      1 äggdonation
      1 Äggdonation
     24 äggen
     15 Äggen
     40 ägget
      5 Ägget
      3 äggets
      1 äggfollikler
      1 äggformade
      1 Äggkläckningen
      1 äggkläckningsmaskin
      1 äggkokonger
      2 äggläggning
      2 äggläggningen
      5 äggledare
      7 äggledaren
      3 äggledarinflammation
      8 äggledarna
      1 Äggledarna
      1 agglomererar
     14 ägglossning
      1 Ägglossning
      2 ägglossningar
     26 ägglossningen
      2 Ägglossningen
      1 ägglossningscykler
      1 ägglossningstest
      1 agglutinationtpha
      1 äggmök
      1 äggproducenten
      2 aggregat
      3 aggregatet
      6 aggression
      3 aggressionen
      3 aggressioner
      1 aggressionsutbrott
     17 aggressiv
     11 aggressiva
      1 aggressivare
     10 aggressivitet
     10 aggressivt
      1 aggreverande
      2 äggrund
      5 äggrunda
      2 äggskal
      2 äggskalet
      1 äggskalsförtunning
      3 äggstock
      1 Äggstock
     18 äggstockar
      1 Äggstockar
     24 äggstockarna
      7 Äggstockarna
      3 äggstockarnas
      5 äggstocken
      9 äggstockscancer
      3 Äggstockscancer
      1 äggstockscystor
      1 äggstocksinflammation
      1 äggstockssnitt
      1 äggstockssvulst
      1 äggtand
      1 äggulan
      4 äggvita
      1 äggvitan
      1 agi
      7 agitation
      2 agiterade
      3 agkistrodon
      7 ägna
      1 ägnad
      5 ägnade
     19 ägnar
      3 ägnas
      1 ägnat
      1 agneta
      1 agnetha
      1 agno
      4 agnosi
      1 agnosia
      1 agnostiker
      1 ägo
      3 ägodelar
      3 agonism
      2 agonist
      2 agonister
      1 agonistes
      1 agora
     20 agorafobi
      1 agorafobiker
      1 agorafobiska
      1 agrafe
      4 agraff
      1 agraffer
      1 agraffspänne
      1 agrammatism
      2 agranulocytos
      1 agria
      2 agrobacterium
      1 agrostemma
      4 ägs
      8 ägt
      1 ahfpreparat
      1 ahitofel
      1 ahlbergs
      1 ahlberts
      4 ahn
      1 ahvaz
      1 aia
      1 aid
     45 aids
      1 aidsdefinierande
      1 aidsepedimin
      1 aidsepidemin
      3 aidsfallet
      1 aidsforskningen
      1 aidskommissionen
      2 aidspatienter
      1 aidsprevention
      1 aidsrelaterad
      2 aidsrelaterade
      1 aidssjuk
      1 aidwa
      1 aifa
      1 aijing
      1 aikido
      1 aikidoinstruktör
      1 aikidons
      2 aina
      1 ainfektion
      3 ainsworth
      1 ainufolket
      2 aip
      2 air
      1 airtruk
      5 airway
      1 aisth�sis
      3 a�j
      1 ajax
      1 ajcc
      1 ajovanolja
     12 åka
      1 akaciablad
      2 akademi
      2 akademien
      1 akademiens
      2 akademiker
      1 akademikerförbundet
      1 akademinska
     17 akademisk
     14 akademiska
      4 akademiskt
      1 akalkyli
      1 akasha
      1 akatesier
      7 akatisi
      1 akedia
      1 akema
      8 åker
      1 åkerjordarna
      1 åkerklätt
      2 Åkerklätt
      3 åkermark
      1 Åkermarken
      1 åkermarkskalkning
      1 åkerogräs
      1 Åkerrök
      1 Åkesson
      1 akillessenan
      1 akinesi
      3 akinetisk
      4 akk
      3 åklagare
      1 Åklagaren
      2 åklagarmyndighet
      1 aklorhydri
     10 akne
      1 akneliknande
     17 åkomma
     13 åkomman
      4 Åkomman
      1 åkommans
     27 åkommor
      4 Åkommor
      9 akondroplasi
      1 akonitin
      1 akrani
      4 åkrar
      2 akrokordon
      1 akrolein
     57 akromegali
      4 akromegalin
      2 akromegaloid
      1 akromegaloidism
      4 akronym
      1 akronymen
      2 akrosom
      5 akrosomen
      1 akrylamid
      1 akrylat
      1 akrylater
      1 akrylatplast
      1 akrylfiber
      1 akrylplast
      1 åksjuk
      2 åksjuka
      1 Åksjuka
      1 åksjukebesvär
      1 akt
     21 äkta
      2 Äkta
      1 aktar
      1 åkte
      7 äktenskap
      9 äktenskapet
      1 äktenskapliga
      5 äktenskapsbrott
      1 äktenskapshinder
      1 äktenskapslöfte
      1 äktenskapsskillnad
      1 akter
      1 äkthet
      1 aktiebolag
      1 aktiemarknaden
      6 aktier
      1 aktinfilament
      3 aktiniderna
      2 aktinobakterier
      1 aktinoiderna
      5 aktinolit
      1 aktinomyceter
      3 aktinos
      2 aktioner
      1 aktionoliten
      1 aktionsinriktat
      9 aktionspotential
      2 aktionspotentialen
      1 aktionspotentialens
      2 aktionspotentialer
      1 aktis
     70 aktiv
     64 aktiva
      2 aktivator
     11 aktivera
      5 aktiverad
      4 aktiverade
      1 aktiverades
      2 aktiverande
     23 aktiverar
     57 aktiveras
      4 aktiverat
     30 aktivering
      6 aktiveringen
      1 aktiveringssignal
      1 aktiveringssystemet
      1 aktivister
     98 aktivitet
     48 aktiviteten
     58 aktiviteter
      5 aktiviteterna
      1 aktivitetsanalys
      2 aktivitetsanalysen
      3 aktivitetsförmåga
      1 aktivitetsförmågan
      2 aktivitetsgrad
      1 aktivitetsmönster
      2 aktivitetsträning
      1 aktivitetsutförande
      7 aktivitetsvetenskap
      1 aktivitetsvetenskapen
      2 aktivitetsvetenskapens
      1 aktivitetsvetenskapsprogrammet
      2 aktivslamprocess
      3 aktivslamprocessen
     38 aktivt
      1 aktör
     11 aktörer
      3 aktörerna
      1 aktualiserar
     13 aktuell
     30 aktuella
     22 aktuellt
      1 aktuta
      2 akupressur
      1 akupukturen
      1 akupunktörer
     23 akupunktur
      1 akupunkturanvändning
      1 akupunkturbehandling
      3 akupunkturens
      1 akupunkturkongressen
      2 akupunkturmetoder
      1 akupunkturnålar
      1 akupunkturpunkter
      1 akupunkturpunkterna
      1 akurvan
      2 akustik
      1 akustikbyrån
      2 akustiker
      1 akustikfirmorna
      2 akustikkonsult
      1 akustikkonsulten
      2 akustikusneurinom
      8 akustiska
      1 akustiskt
    189 akut
     69 akuta
      1 akutavdelningar
      2 akuten
      1 akutfall
      1 akutfasprotein
      1 akutfasproteiner
      1 akutfasreaktanter
      1 akutkirurgisk
     11 akutläkare
      1 akutläkaren
      1 akutläkemedel
      3 akutmottagning
      2 akutmottagningar
      8 akutmottagningen
      1 akutmottagnings
      1 akutomedelbar
      2 akutppiller
      2 akutppillret
      1 akutprov
      2 akutsjukhus
      4 akutsjukvård
      1 akutsjukvården
      1 akutsjukvårdsspecialiteten
      2 akutskedet
      1 akutspruta
      2 akuttestet
      1 akuttillstånd
      2 akutvård
      1 akutvårdsavdelning
      1 akutverksamheten
      1 akvamarin
      1 akvariefiskar
      1 akvarium
      3 akvatiska
      1 akzo
     32 al
     10 ala
      2 alabama
      1 ålagda
      2 ålägga
      2 ålägger
      5 alan
      3 Åland
      2 alanin
      2 alaninaminotransferas
      2 alarm
      1 alarmämnen
      2 alarmferomoner
      1 alarmreaktion
      1 alarmsignaler
      2 alaska
      9 alat
      1 alatvärden
      5 alba
      1 albaner
      3 albendazol
     21 albert
      1 alberta
      1 albertus
      2 albicans
      3 albina
     21 albinism
      1 albinismen
      1 albinistiska
      2 albinistiskt
      3 albino
      1 albinodjur
      1 albinofärgad
      1 albinofärgerna
      1 albinoteckning
      1 albinsim
      2 albopictus
      1 albrecht
      1 albrekt
      1 albuginea
      1 album
      2 albumen
      2 albumet
     11 albumin
      1 albuminproduktion
      1 alby
      1 albysjöns
      1 alcohol
      2 alcoholism
      1 alcoholismus
      1 alcor
      1 ald
      1 aldara
      1 alddrabbade
      1 aldehyd
      2 aldehyder
      1 aldehydgrupp
    261 ålder
      1 Ålder
      4 ålderdom
      1 Ålderdom
      6 ålderdomen
      2 ålderdomens
      2 ålderdomlig
      2 ålderdomligt
      1 ålderdomshem
      1 ålderdomssvaghet
      1 ålderdomstecken
      1 åldergruppen
      1 Åldermässigt
     26 åldern
      3 Åldern
      1 åldersangivelsen
      1 åldersberoende
      1 åldersbestämma
      1 åldersbestämning
      1 åldersbetingad
      2 åldersdiabetes
      1 åldersdiabetesinsulinoberoende
      1 åldersfläckar
      2 åldersförändring
      1 åldersgräns
      5 åldersgrupp
      6 åldersgruppen
      8 åldersgrupper
      1 åldersgrupps
      1 åldersintervall
      2 åldersintervallet
      1 ålderskategorier
      1 ålderskrämpor
      1 Åldersmässigt
      1 ålderspåverkan
      1 åldersperiod
      2 åldersrelaterad
      6 åldersrelaterade
      1 åldersrelaterat
      1 åldersstandardiserad
      1 åldersstrukturerad
      1 ålderssvaghet
      1 ålderssymtom
      1 ålderssynt
      3 ålderssynthet
      1 Åldersuppskattningarna
      1 åldersutredning
      1 åldersvariationer
      1 åldersynthet
      1 aldh
      1 aldomet
      1 aldoncia
      2 aldosteron
      2 aldosteronism
      1 åldrade
     26 åldrande
      3 Åldrande
      1 åldrandeprocessen
      7 åldrandet
      3 åldrandets
     28 åldrar
     14 åldrarna
      7 åldras
    237 äldre
     21 Äldre
      3 äldreboende
      1 äldreboenden
      5 äldreomsorg
      1 Äldreomsorg
      3 äldreomsorgen
      1 äldrepolitik
      1 äldres
      2 äldrevård
     93 aldrig
      1 åldringar
      1 Åldringar
      1 åldringslinjer
      1 åldringsprocessen
      3 äldst
     37 äldsta
      1 alec
      1 alejandro
      1 aleksej
      1 alerta
      1 alerthet
      3 alessandro
      7 alexander
      1 alexandergradering
      3 alexandertekniken
      1 alexandre
      9 alexi
      3 alexier
      1 alexin
      1 alexithymia
     12 alexitymi
      1 alf
      7 alfa
      1 alfaantitrypsin
      2 alfaantitrypsinbrist
      1 alfaantitrypsinnivån
      1 alfabåren
      1 alfabeten
      4 alfabetet
      2 alfabetisk
      1 alfabindingar
      1 alfabindningar
      2 alfabindningarna
      1 alfafetoprotein
      1 alfaglukos
      1 alfaglukosidashämmare
      1 alfaglykosidbindning
      1 alfaglykosidbindningar
      1 alfahelixar
      3 alfahemolytiska
      1 alfahydroöstron
      1 alfahydroxyöstron
      1 alfaintegriner
      2 alfametyldopa
      1 alfametylnoradrenalin
      1 alfamotorneuron
      1 alfaöstron
      2 alfapartiklar
      1 alfareceptorblockerare
      1 alfareceptorer
      1 alfastrålande
      3 alfastrålning
      1 alfastrålningen
      1 alfastreptokocker
      1 alfasynuklein
      2 alfavirus
      7 alfred
      1 alfredsson
      1 alfvén
      5 älg
      1 algdödande
      1 älgens
     10 alger
      1 algeriet
      1 Älgfluga
      1 Älgflugan
      1 älgflugor
      1 algicid
      1 älglus
      1 algologi
      1 algoritmer
      2 algos
      2 ali
      1 aliberts
      2 alice
      1 alien
      1 alienum
      1 alifatisk
      1 alifatiskt
      2 åligger
      1 aliknande
      1 alimentarius
      1 alimlouis
      1 aliskiren
      1 alive
      1 alizarin
      1 alkali
      1 alkaliejodider
      2 alkalier
      2 alkalimetaller
      1 alkalina
      1 alkaliserade
      2 alkalisk
      6 alkaliska
      2 alkaliskt
      1 alkaloid
      6 alkaloiden
      7 alkaloider
      3 alkaloiderna
     15 alkalos
      1 alkalosen
      1 alkan
      2 alkaseltzer
      1 alkemi
      1 alkemilitteratur
      1 alkemins
      1 alkemist
      4 alkemister
      1 alken
      2 alkener
    118 alkohol
      7 alkoholabstinens
      1 alkoholabstinenssyndromet
      2 alkoholbaserade
      1 alkoholbaserat
      7 alkoholberoende
      1 alkoholberoendet
      2 alkoholbruk
      1 alkoholbrukare
      1 alkoholcirros
      3 alkoholdehydrogenas
      2 alkoholdelirium
      1 alkoholdryck
      5 alkoholdrycker
     10 alkoholen
      1 alkoholens
     36 alkoholer
      2 alkoholerna
      1 alkoholextrakt
      1 alkoholförbudet
      2 alkoholförgiftning
      1 alkoholförgiftningens
      1 alkoholforskare
      2 alkoholförtäring
      1 alkoholfria
      1 alkoholgeler
      1 alkoholgruppen
      2 alkoholhalt
      1 alkoholhalten
      6 alkoholhaltiga
      1 alkoholhepatit
      5 alkoholintag
      1 alkoholintaget
     17 alkoholism
      2 alkoholismen
      1 alkoholismens
      2 alkoholist
      7 alkoholister
      1 alkoholisters
      1 alkoholkoncentrationen
      7 alkoholkonsumtion
      1 alkoholkonsumtionen
      1 alkoholleverskada
      1 alkohollösning
     11 alkoholmissbruk
      1 alkoholmissbruket
      1 alkoholmolekylerna
      1 alkoholöverkonsumtion
      1 alkoholparanoia
      1 alkoholpåverkade
      3 alkoholpåverkan
      1 alkoholpåverkat
      1 alkoholproblem
      2 alkoholrelaterade
      2 alkoholrus
      1 alkohols
      1 alkoholskatt
      1 alkoholsyndrom
      1 alkoholtillförseln
      2 alkoholutlöst
      2 alkoholutlösta
      1 alkometer
      1 alkyldimetylbensylammoniumklorid
      1 alkylerande
      1 alkylering
      2 alkyner
     88 all
    789 alla
      1 allah
      1 allander
      1 allanmcormack
      1 alldagliga
      1 alldagligt
     11 alldeles
      3 allehanda
      1 allelen
      4 alleler
      2 allelerna
      1 allelopati
      1 allelopatiska
      1 allenarådande
      1 allergan
     27 allergen
      2 allergena
      2 allergenen
      5 allergener
      2 allergenerna
      2 allergenet
      2 allergenextrakt
      1 allergenextrakten
      1 allergenkälla
      1 allergens
      1 allergenstandardisering
      1 allergent
     58 allergi
      1 allergiåtgärdsplan
      5 allergichock
      1 allergidiagnos
      1 allergidiagnostiken
     14 allergier
     14 allergiframkallande
      2 allergiker
      1 allergikerna
      3 allergiliknande
      1 allergimediciner
      4 allergin
      1 allergireaktion
     41 allergisk
     47 allergiska
      4 allergiskt
      1 allergisprutor
      2 allergisyndromet
      1 allergitestade
      4 allergitester
      3 allergiutredning
      1 allergivaccinering
      1 allergologi
      1 allesammans
      1 allgemeinbildung
      1 allgemeinmedizin
      1 alliance
      4 allicin
      1 alliera
      3 allierade
      1 allierades
      1 allierat
      1 alligatorer
      1 allindia
      1 allm
     60 allmän
      1 allmänbildad
      4 allmänbildning
      1 allmänbildningsnivå
      7 allmänfarlig
      4 allmänfarliga
      3 allmängiltiga
      2 allmängods
      1 allmänhälsa
      1 allmänhänseende
     77 allmänhet
     15 allmänheten
      1 allmänhetens
      1 allmänhygienen
      1 allmäninfektioner
      1 allmänkirurger
      1 allmänkirurgin
      5 allmänläkare
      1 allmänläkaresköterskor
      1 allmänläkarkompetens
      1 allmänljus
      1 allmänmänsklig
      1 allmänmänskliga
     11 allmänmedicin
      3 allmänmedicinare
      2 allmänmedicinaren
      1 allmänmedicinen
      1 allmänmedicinska
      1 allmänn
     70 allmänna
      1 allmänpåverkan
      1 allmänpsykiatrin
      1 allmänreaktioner
      1 allmänsjukdom
      2 allmänsymptom
      1 allmänsymtom
     76 allmänt
      1 allmäntandläkare
      1 allmäntandvården
      7 allmäntillstånd
      7 allmäntillståndet
      1 allmäntjänstgöring
      1 allmoge
      3 allmogen
      1 allmosor
      1 alloderm
      3 allodyni
      1 allogen
      1 allomon
      1 allopurinol
      1 allostas
      1 alloster
      1 allostera
      1 allotropa
      1 allotropi
      2 allotropiska
      1 allotropiskt
     58 allra
     54 alls
      1 allsidig
      1 allsmäktiga
    391 allt
      5 allteftersom
      1 alltereftersom
      1 alltfler
     49 alltför
    217 alltid
      7 alltifrån
      1 allting
      6 alltjämt
     16 alltmer
    219 alltså
      3 alltsedan
      1 allusionen
      1 allvaligare
     10 allvar
      1 allvaret
    115 allvarlig
    156 allvarliga
     39 allvarligare
      1 allvarligast
     16 allvarligaste
      2 allvarlighet
      4 allvarlighetsgrad
      7 allvarlighetsgraden
     57 allvarligt
      2 allvetande
      1 allylalkohol
      1 allylamin
      1 allylisotiocyanat
      4 allylklorid
      1 allylkloridförgiftning
      1 allylsilan
      1 allylsulfensyra
      1 allyn
      1 almajidrefref
      2 almanackor
      2 almansur
      1 almindelig
      1 alnarp
      1 alo
      4 aloe
      1 aloh
      1 alois
      1 alooh
      2 alopecia
      3 alperna
      1 alpestris
      2 alpgullregn
      1 alpgullregnets
      1 alpha
      1 alphametylfenetylamin
      2 alpinum
      2 alprazolam
      1 alpstegring
      1 alpstormhatt
      1 alpstormhatten
      1 alptopparna
      1 alqasim
      1 alrazi
      4 alruna
      5 alrunan
      3 alrunans
      2 alrunorna
      2 als
      2 älska
      1 älskade
      1 älskande
      1 älskar
      1 älskare
      1 älskarinnors
      1 älskat
      1 älsklig
      7 alstra
      5 alstrar
      6 alstras
      3 alt
      1 ältande
      1 alteplas
      2 alternaria
     94 alternativ
     38 alternativa
      4 alternativen
      7 alternativet
      1 alternativkomplement
     14 alternativmedicin
     10 alternativmedicinen
      8 alternativmedicinsk
     10 alternativmedicinska
      1 alternativmedicinskt
      2 alternativnamn
     52 alternativt
      1 alternativvården
      1 alternera
      1 alternering
      2 altitud
      2 altitude
      1 altituden
      1 altman
      2 altruism
      1 alumini
     17 aluminium
      2 aluminiumbaserade
      1 aluminiumet
      1 aluminiumhalter
      5 aluminiumhydroxid
      1 aluminiumhydroxiden
      1 aluminiumjoner
      3 aluminiumklorid
      2 aluminiumkloridhydrat
      3 aluminiumoxid
      1 aluminiumoxidhydroxid
      1 aluminiumsalt
      1 aluminiumsalter
      1 aluminiumsalterna
      1 aluminiumupptagning
      2 aluminiumzirkonium
      1 alumni
     10 alun
      1 alunbad
      1 alunhaltiga
      1 alunskiffer
      1 alunstift
      1 alva
      1 alvar
      2 alvarezi
      1 alvarligt
      2 alvastra
      2 alvedon
      1 alveol
      6 alveolär
      3 alveolära
      1 alveolarkapillärerna
      5 alveolen
      7 alveoler
     17 alveolerna
      1 alveoli
      2 alveolit
      1 alveolkapillärväggen
      1 alveolväggarna
      1 alversta
      1 alvesta
      1 alvestaepidemin
      1 alvin
      1 älvor
      1 älvors
      1 alzahrawi
      3 alzheimer
      2 alzheimerpatienter
     22 alzheimers
      1 alzheimerssymptom
      4 am
      1 ama
      1 amadeus
      1 amae
      4 amalgam
      1 amalgamer
      1 amalgamförgiftning
      1 amalgamfyllningar
      1 amalgamsanering
      1 amalgamspån
      1 amalgamutborrning
      2 amandiana
      1 amanita
      1 amanitaceae
      2 amanitin
      3 amantadin
      1 amarae
      1 amaranth
      1 amaranthus
      1 amaris
      1 amaroneviner
      1 amartya
      2 amaryllisväxter
      1 amatörer
      1 ämbete
      2 ämbeten
      1 ämbetsmän
      1 ambition
      2 ambitionen
      1 ambitionerna
      1 ambitiösa
      1 ambivalens
      1 amblycera
      1 ambrahamitiska
      2 ambroise
      1 ambros
      1 ambrotyper
      1 ambulance
      8 ambulans
      1 ambulansbårar
      1 ambulansbilar
      2 ambulansen
      1 ambulanser
      1 ambulansfordon
      4 ambulanspersonal
      3 ambulanssjukvård
      3 ambulanssjukvårdare
      1 ambulanssjukvårdaren
      2 ambulanssjukvården
      1 ambulare
      1 ambystoma
      2 ambystomatidae
      3 amenorré
      3 america
     20 american
      1 americana
      1 americatävling
      2 americium
     21 amerika
      1 amerikan
      6 amerikanen
      3 amerikaner
      2 amerikanerna
     13 amerikansk
     62 amerikanska
      4 amerikanskan
     16 amerikanske
      6 amerikanskt
      2 amerikas
      1 amerikavinnare
     46 amfetamin
      1 amfetaminalkaloid
      2 amfetaminberoende
      1 amfetaminberoendet
      1 amfetaminberoendets
      1 amfetaminbrukaren
      1 amfetaminchchchnhch
      2 amfetaminderivat
      1 amfetaminepidemins
      1 amfetaminer
      3 amfetaminet
      4 amfetaminets
      1 amfetaminfribasen
      3 amfetamingruppen
      1 amfetaminhydroklorid
      1 amfetaministen
      3 amfetaminliknande
      5 amfetaminmissbruk
      3 amfetaminmissbrukare
      1 amfetaminmissbruket
      2 amfetaminmolekylen
      1 amfetaminpåverkade
      1 amfetaminpåverkades
      1 amfetaminpåverkan
      1 amfetaminpreparaten
      1 amfetaminpsykosen
      2 amfetamins
      5 amfetaminsalt
      2 amfetaminsalter
      2 amfetaminsulfat
      1 amfetamintabletter
      2 amfibol
      1 amfibola
      6 amfiboler
      1 amfibolernas
      1 amfibolgrupper
      1 amfibolit
      1 amfibolmineral
      1 amfibolos
      1 amfolyt
      2 amfotericin
      1 amination
      9 amineptin
      1 amineptinmolekylen
      6 aminer
      1 aminfluorid
      1 amingrupp
      1 amingrupper
      1 åminnelse
      1 aminofenol
      1 aminoglykosid
      2 aminoglykosider
      1 aminogrupp
      1 aminohydroxifenyl
      1 aminokvävet
      1 aminolevulinat
      3 aminolevulinsyra
      1 aminooxopentansyra
      3 aminosalicylsyra
      6 aminosyra
      6 aminosyran
      1 aminosyrasekvensen
      1 aminosyrebärare
     28 aminosyror
      3 aminosyrorna
      1 aminoterminalt
      1 aminotransferaser
      1 aminotransferasstegring
      1 aminoxidas
      1 amiodaron
      2 amitokondriska
      1 amitriptylin
      2 amitrol
      1 aml
      8 amma
      3 ammande
      2 ammar
      2 ammas
      1 ammats
     29 ammoniak
      3 ammoniaken
      1 ammoniakframställningen
      1 ammoniakhalten
      1 ammoniaklösning
      1 ammoniaksilverlösningar
      1 ammoniakutsläpp
      2 ammonium
      1 ammoniumförening
      2 ammoniumhydroxid
      1 ammoniumjonen
      2 ammoniumjoner
      1 ammoniumkatjon
      1 ammoniumnitrat
      1 ammoniumperteknat
      3 ammunition
      1 ammunitionvapen
      1 amn
      2 ämnad
      1 amnade
      2 ämnade
     87 ämne
    203 ämnen
      7 Ämnen
     17 ämnena
      3 ämnens
      5 ämnes
      2 ämnesbeteckning
      7 amnesi
      1 amnesia
      1 ämnesinnehåll
      1 amnesisyndrom
      2 ämnesklassen
      1 ämnesområde
      2 ämnesområden
      1 Ämnesområden
      1 ämnesområdena
      4 ämnesområdet
      2 Ämnesområdet
     21 ämnesomsättning
      1 Ämnesomsättning
     12 ämnesomsättningen
      2 Ämnesomsättningen
      2 ämnesomsättningshormoner
      2 ämnesomsättningshormonerna
      3 ämnesomsättningsrubbningar
      1 ämnesomsättningssjukdom
      3 ämnesomsättningssjukdomar
      1 Ämnesomsättningssjukdomar
      1 ämnesrubriker
      1 Ämnesrubrikerna
      1 ämnesspecifika
      1 amnesti
    110 ämnet
     65 Ämnet
      5 ämnets
      4 Ämnets
     20 amning
      1 amningar
      2 amningarna
      6 amningen
      1 amningens
      1 amningshormoner
      1 amningsnapp
      1 amningspsykos
      1 amningsställning
      1 amningsteknik
      1 amningstiden
      3 amnionvätskan
      3 amöbadysenteri
      1 amöbaorsakad
      8 amöbor
      2 amöborna
      4 amok
      1 amon
      1 amorbåge
      2 amorf
      2 amosit
      1 amotio
      5 amoxicillin
      1 ampa
      1 ampareceptorn
      1 ampelskära
      3 ampere
      3 amperemeter
      2 amperemetern
      1 amperemetrar
      1 amphicarpos
      1 amphotericin
      3 ampicillin
      1 amplifiera
      1 amplifieringar
      6 amplitud
      1 amplituden
      1 amplitudmodulerad
      1 amplitudvariation
      2 amp�re
      3 amps
      2 ampull
      1 ampulla
      1 ampullen
      6 amputation
      1 amputationer
      2 amputera
      1 amputerade
      1 amputerades
      1 amputeras
      1 amputerat
      4 ams
      3 amsterdam
      1 amulett
      1 amuletten
      2 amusi
     17 amygdala
      1 amygdalae
      7 amygdalin
     10 amylas
      1 amylaser
      1 amylaserna
      4 amyloid
      1 amyloida
      1 amyloidernas
      4 amyloidos
      2 amyloidoser
      1 amylopektin
      1 amylos
      1 amylovora
      1 amylum
     10 an
   1112 än
      5 Än
      6 ana
      2 anaanhängare
      2 anabol
     16 anabola
      1 anabolt
      1 anacardiaceae
      5 anaerob
     18 anaeroba
      3 anaerobt
      1 anaesthetics
      1 anafranil
     12 anafylaktisk
      2 anafylaktiska
      1 anafylaktoida
     76 anafylaxi
      1 anafylaxibehandling
      1 anafylaxifallen
      1 anafylaxin
      2 anagyroides
      1 anakulturen
      4 anal
      5 anala
      1 analens
      1 analfissur
      8 analgetika
      2 analgetikum
      1 analgetiska
      3 analkanalen
      3 analkuddar
      3 analkuddarna
      7 analog
     12 analoga
      1 analogdigitalomvandlare
      5 analogi
      1 analogier
      2 analogin
      6 analogt
      2 analöppning
     12 analöppningen
      1 analpapiller
      1 analpropp
      1 analsäcksinflammation
      5 analsex
      1 analsfinktern
      1 analsfinkterns
      4 analt
      1 analtampong
     33 analys
      2 analysatorer
      1 analysautomat
      1 analysautomater
      7 analysen
      1 analysens
     12 analyser
     15 analysera
      4 analyserade
      4 analyserar
      6 analyseras
      1 analyserats
      2 analyserna
      1 analysinstrument
      4 analysis
      1 analysmedel
      3 analysmetoder
      1 analyssis
      3 analyst
      2 analysverktyg
      1 analyten
      3 analytiker
      1 analytikern
      2 analytisk
      1 analytiska
      1 analytiskt
      1 anammar
      1 anammat
      9 anamnes
      1 anamnesbaserad
      4 anamnesen
      1 anamnesis
      1 anamorph
      1 ananas
      1 anaplasma
      1 anaplasmabakterien
      1 anaplasmainfektionen
      3 anaplastisk
      1 anarkister
      1 anarkistfilosofen
      1 anarkokapitalism
      1 anasarka
      2 anastomos
      2 anastomoser
      2 anastomoserande
      1 anastrozol
      1 anatma
      1 anatoli
      1 anatom
      1 anatomen
     27 anatomi
      1 anatomibok
      4 anatomin
      8 anatomisk
     18 anatomiska
      6 anatomiskt
      1 anatoxin
      1 anatripsisven
      1 anatta
      2 anaxagoras
      1 anbragta
      1 anbringade
      4 anbringas
      1 anbringats
     93 and
      1 änd
      2 anda
     40 ända
      6 Ända
     78 ändå
      1 Ändå
     33 ändamål
      1 Ändamål
      7 ändamålet
      2 Ändamålet
      2 ändamålsenlig
      3 ändamålsenligt
      1 ändamålslösa
      9 andan
      4 ändan
      1 andante
     14 andar
      4 ändar
      1 andare
      1 andarkrafterförfäder
      3 andarna
      2 ändarna
      1 andarnaförfäderna
      1 andarnas
     92 andas
      1 andats
      1 ändavslut
      1 anddr
     22 ande
      8 ände
      1 andedop
     20 andedräkt
      3 andedräkten
      1 andedrömvärlden
      1 andegåvor
     54 andel
     62 andelen
      1 Ändelsen
      1 andelsrekommendation
      1 andemagiker
     12 anden
     20 änden
      4 andens
      1 anderna
     11 anders
      1 andersensaga
      1 andersonfabrys
      2 andersson
      4 anderstorp
      1 andesit
      1 andestoff
     18 andetag
      2 andetagen
      1 andetaget
      1 andetagminut
      2 andetagsfrekvensen
      1 andeutdrivning
      3 andevärlden
      1 andevärldendrömvärlden
      1 andeväsen
     10 andfåddhet
      1 andfåglar
      1 andingsmask
     14 andlig
     16 andliga
      3 andlighet
      1 andligt
      1 andligtexistentiellt
      1 andligtmentala
      1 ändlös
      1 ändmål
     49 andning
     30 andningen
      3 andningens
      2 andnings
      2 andningsapparat
      2 andningsapparaten
      1 andningsballong
      1 andningsballonger
      1 andningsbesvär
      1 andningscentra
      4 andningscentrum
      4 andningsdepression
      1 andningsdepressionen
      1 andningsdepressiva
      1 andningsförlamning
      1 andningsförmåga
     12 andningsfrekvens
      6 andningsfrekvensen
      4 andningsgas
      1 andningsgymnastik
      1 andningshinder
      1 andningshjälp
      2 andningskontroll
      1 andningsljud
      2 andningsljuden
      1 andningsluften
      1 andningsmönstret
      1 andningsmuskler
      1 andningsmusklerna
      4 andningsmuskulaturen
      1 andningsneuron
      2 andningsöppning
      3 andningsorgan
      4 andningsorganen
      1 andningsorgansfel
      2 andningsövningar
      1 andningspassagen
      4 andningsproblem
      1 andningsproblemet
      1 andningsreflexen
      2 andningsreglerande
      1 andningsregleringen
      1 andningsrelaterad
      1 andningsrör
      2 andningsrörelser
      1 andningsröret
      2 andningsrytm
      3 andningsrytmen
      1 andningssgasens
      1 andningssignaler
      2 andningsskydd
      7 andningsstillestånd
      1 andningsstödsproblem
      1 andningsstörningar
      3 andningsstörningarna
      1 andningsstörningsepisoder
      9 andningssvårigheter
      1 andningssvårigheterna
      2 andningssvikt
      3 andningssystemet
      1 andningstakt
      2 andningsteknik
      1 andningstekniker
      7 andningsuppehåll
      1 andningsuppehållen
      1 andningsuppehållens
      4 andningsvägar
     12 andningsvägarna
      1 andningsvägen
      1 andningsvolymen
     17 andnöd
      1 andnor
      1 ändöglor
      1 andosteron
      1 ändplatta
      1 ändplattor
      1 ändpunkter
   1941 andra
     23 ändra
      5 ändrad
      6 ändrade
      1 Ändrade
     14 ändrades
      1 andradivisionen
     21 ändrar
      1 ändrarna
     22 andras
     18 ändras
      8 ändrat
      7 ändrats
     17 andre
      2 andré
      1 andrea
      2 andreas
      1 andrémarie
      5 andres
      3 andrew
      4 ändring
      2 Ändring
      6 ändringar
      1 Ändringar
      1 ändringarna
      2 androblastom
      1 androcymbium
      8 androgena
      1 androgenen
     27 androgener
      7 androgenerna
      1 androgenernas
      4 androgenokänslighet
      1 androgenokänslighetssyndrom
      3 androgenreceptorn
      1 androgenvärden
      1 androlog
      1 androloger
      1 andrologi
      1 andrologin
      2 andromachus
      3 andropaus
     17 androstendion
      1 androstendionen
      1 andry
      1 andtäppa
      2 ändtarm
     22 ändtarmen
      3 Ändtarmen
      2 ändtarmens
      1 ändtarmscancer
      1 ändtarmsöppning
      3 ändtarmsöppningen
      1 ändtarmssköljning
      1 ändtarsmöppningen
      1 andy
      1 anell
     29 anemi
      1 anemier
      1 anemisk
      4 anemone
      1 anemoner
      5 anencefali
      2 anencefaliska
      1 anencefalt
      1 anencephali
      1 anenue
      1 anervan
     24 anestesi
      1 anestesigas
      1 anestesigasen
      1 anestesiläkaren
      1 anestesiläkemedel
      1 anestesimedel
      3 anestesin
      1 anestesins
      3 anestesiolog
      1 anestesiologer
      3 anestesiologi
      1 anestesiologin
      1 anestesiologisk
      2 anestesipersonal
      2 anestetika
      3 anestetikum
      1 anestetiska
      1 anetolhalten
      1 aneuploida
      2 aneuploidi
     11 aneurysm
      3 aneurysma
      1 aneurysmbildning
      1 aneurysmen
      1 aneurysmer
      1 aneurysmet
     58 anfall
      2 anfalla
      1 anfallande
      4 anfallen
      4 anfaller
      6 anfallet
      1 anfallna
      4 anfallsfria
      3 anfallsfrihet
      1 anfallstyper
      1 anfallsutlösande
      1 anfallsvis
      1 anförare
      1 anförd
      1 anförde
      1 anfördes
      1 anförtro
      1 anförtrodd
      1 anförts
      9 ånga
     14 angående
      1 ångan
      3 ängar
      2 angår
      6 angav
      4 angavs
      1 ångbad
      1 Ångbad
      2 ångbastu
      9 ange
      2 angeion
      2 ängel
      2 angelägenhet
      2 angelägenheter
      2 angeläget
      3 angeles
      1 angelesolympiaden
      1 angelo
      1 angelologi
      1 ängen
      1 angenäma
      1 angenämt
     43 anger
      5 ånger
      1 ångerkänslor
      1 Ångermanälvens
     64 anges
      2 ångesstörningar
     94 ångest
      5 Ångest
      1 ångestattack
      1 Ångestattacken
      7 ångestdämpande
      1 ångestdrivande
     17 ångesten
      1 Ångesten
      1 ångestframkallande
      1 ångestfri
      1 ångestfylld
      2 ångestfyllda
      1 ångestfyllt
      2 ångestkänslor
      2 ångestkänslorna
      1 ångestlindrande
      1 Ångestlindrande
      1 ångestlindring
      1 ångestminskning
      2 ångestnivå
      2 ångestnivån
      1 ångestreaktioner
      1 Ångestreaktioner
      1 ångestreduktion
      1 ångestrelaterade
      1 ångestsjukdomar
      1 ångestskapande
      6 ångeststörning
     18 ångeststörningar
      4 Ångeststörningar
      1 ångeststörningarnas
     13 ångestsyndrom
      1 Ångestsyndrom
      1 ångestsystem
      5 ångesttillstånd
      1 ångestupplevelser
      1 ångestutlöst
      1 ångestväckande
      3 angett
      1 angetts
      2 ångform
      1 angigenes
      3 angina
     10 angiogenes
      1 angiogenesen
      4 angiogeneshämmare
      7 angiografi
      1 angiografiskt
      1 angiogram
      1 angiokärl
      1 angiolipom
      4 angiom
      1 angioma
      1 angiomyolipom
      8 angioödem
      1 angioödemet
      1 angioosteohypertrofiskt
      3 angioplastik
      3 angiosarkom
      1 angiospermer
      3 angiospermerna
      1 angiostrongylus
     22 angiotensin
      1 angiotensine
      3 angiotensinkonverterande
      3 angiotensinogen
      1 angiotensinogenet
      1 angiotensinreceptorhämmarna
      1 angiotensinreceptorn
      2 angiper
      1 angivelse
      2 angiven
      1 angivet
      2 angivit
      1 angivits
      3 angivna
      1 ångkoka
      2 ångkokning
      1 Ångkokning
      1 änglapotta
      2 änglar
      3 ånglok
      1 Ångloket
      2 anglosaxisk
      2 anglosaxiska
      3 ångor
      1 ångorna
      1 ångpannor
      1 Ångpressade
      1 ångra
      1 ångrade
      8 angränsande
      1 ångras
      1 ångrat
      3 angrep
     36 angrepp
      2 angreppen
      4 angreppet
      1 angreppsmetod
      1 angreppspunkter
      1 angreppspunkterna
      2 angreps
     24 angripa
      1 angripare
      1 angriparna
      4 angripas
      2 angripen
     44 angriper
      2 angripet
      5 angripna
      7 angrips
      4 ängslan
      1 ängsliga
      1 ängsligt
      1 ängsmark
      1 ängsmarker
      1 ångstrykjärnet
      1 angularis
      1 angulatus
      1 anhållan
      8 anhängare
      3 anhängarna
     16 anhedoni
      2 anhedonin
      1 anhidrotisk
      2 anhopning
      8 anhörig
     29 anhöriga
      2 anhörigas
      2 anhörigvården
      1 anhydrider
      1 anil
     12 anilin
      1 anilinblått
      1 anilinfärger
      1 anilingrönt
      2 anilinrött
      1 anilinviolett
      2 animal
      1 animalieproducerande
      1 animalier
      1 animalierna
      9 animaliska
      5 animaliskt
      1 animals
      1 animation
      2 anime
      1 animera
      1 animerade
      1 animerar
      1 animeras
      3 animism
      4 aning
      1 aningen
      2 aniridi
      4 anis
      1 anisakiasis
      1 anisogami
      1 anisokori
      1 anisolja
      1 anisum
      3 anjon
      2 anjoner
      1 anka
      3 änka
      3 ankar
      3 ankara
      1 ankarform
      1 ankas
      1 ankel
      1 ankelklonus
      3 ankeln
      1 änkestöt
      2 anklagad
      2 anklagade
      3 anklagades
      2 anklagar
      1 anklagas
      1 anklagats
      2 anklagelser
      3 anklar
      2 anklarna
      1 anknyter
     16 anknytning
      2 anknytningar
      3 anknytningen
      3 anknytningens
      1 anknytningförmåga
      2 anknytningsbeteendet
      1 anknytningsforskningen
      2 anknytningshistoria
      3 anknytningsmönster
      2 anknytningspersonen
      1 anknytningspersoner
      1 anknytningspersonerna
      1 anknytningsproblem
      1 anknytningsprocesser
      1 anknytningsstrategier
      1 anknytningsteori
      4 anknytningsteorin
      1 anknytningsteorins
      2 anknytningsutvecklingen
      1 ankom
      5 ankomst
      1 ankomsten
      1 ankor
      1 änkor
      1 ankskinn
      4 ankyloserande
     22 anlag
      1 anlagd
      1 anlagda
      3 anlagen
     11 anlaget
      2 anlägga
      1 anlägger
      6 anläggning
      4 anläggningar
      1 anläggningarna
      2 anläggningen
      1 anläggningens
      1 anläggningsrubbningar
      4 anläggs
      1 anlags
      4 anlagsbärande
      3 anlagsbärare
      1 anlagsbärarna
      1 anlända
     10 anlände
      1 anlänt
     53 anledning
     17 anledningar
      9 anledningarna
     35 anledningen
      3 anlita
      2 anlitades
      1 anlitar
      4 anlitas
      1 anlitats
      1 anlöpa
      1 anlöps
      1 anm
      7 anmäla
      8 anmälan
      4 anmälas
      6 anmälda
      1 anmälde
      3 anmäldes
      3 anmälningsplikt
      1 anmälningsplikten
     15 anmälningspliktig
      3 anmälningspliktiga
      1 anmälningsskyldighet
      3 anmäls
      3 anmält
      3 anmälts
      5 anmärkning
      1 anmärkningen
      2 anmärkningsvärd
      3 anmärkningsvärda
      2 anmärkningsvärt
      1 anmärkt
      1 anmodan
      1 ann
      5 anna
      1 annales
      1 annals
    399 annan
     10 annans
      9 annanstans
     80 annars
    861 annat
      1 anne
      1 annemarie
      1 annidalin
      1 annihilera
      1 annika
      1 annons
     25 annorlunda
      1 annorstädes
    138 ännu
      5 Ännu
      1 annua
      1 annueller
      1 annulen
      1 annuus
      1 anod
      4 anoden
      1 anoderm
      1 anodmaterialet
      3 anoftalmi
      5 anomalier
      1 anomalies
      1 anomaloskop
      1 anomaloskopet
      1 anomaloskopi
      2 anomaly
      2 anomi
      1 anomisk
      2 anonym
      6 anonyma
      1 anonymous
      1 anonymt
      2 anopheles
      1 anophelesmygga
      2 anophelinae
      3 anoplura
      1 anoplurerna
      1 anor
      1 anordna
      2 anordnade
      2 anordnades
      2 anordnas
     16 anordning
      1 anordningar
      1 anordningen
      2 anorektala
      4 anorektiker
      5 anorexi
     16 anorexia
      1 anorgasmi
      3 anormala
      1 anoskopi
     12 anosmi
      2 anovulation
      2 anoxi
      1 anoxicitet
     17 anpassa
     15 anpassad
     15 anpassade
      1 anpassades
      8 anpassar
      9 anpassas
      8 anpassat
      3 anpassats
     27 anpassning
      1 anpassningar
      1 anpassningen
      1 anpassningmek
      2 anpassningsförmåga
      1 anpassningsreaktionen
      1 anpassningsreaktioner
      1 anpassningsstöd
     17 anpassningsstörning
      4 anpassningsstörningar
      1 anrikades
      2 anrikas
      3 anrikning
     44 ansåg
     65 ansågs
      1 ansamla
      1 ansamlad
      4 ansamlades
      1 ansamlar
     26 ansamlas
      3 ansamlats
     20 ansamling
      4 ansamlingar
      1 ansamlingarna
      3 ansamlingen
      2 ansats
      1 ansatsen
      5 ansatsrör
      6 ansatsröret
      2 ansätter
      1 ansatzrohr
      3 anse
      1 ansedd
      1 ansedda
      3 anseende
      2 ansenlig
     80 anser
    243 anses
      5 ansett
     16 ansetts
     16 ansikte
      1 ansiktebr
      7 ansikten
      1 ansiktena
      1 ansiktes
     53 ansiktet
      1 ansiktets
      1 ansiktigenkänning
      2 ansikts
      1 ansiktsbehandligar
      6 ansiktsblindhet
      1 ansiktsdata
      2 ansiktsdrag
      1 ansiktsdragen
      6 ansiktsförlamning
      1 ansiktsförlamningen
      1 ansiktsformen
      1 ansiktshalvan
      1 ansiktshalvans
      1 ansiktshår
      1 ansiktshud
      1 ansiktsinfektioner
      1 ansiktslyft
      4 ansiktsmask
      1 ansiktsmasker
      1 ansiktsmimiken
      2 ansiktsmuskler
      1 ansiktsmusklerna
      1 ansiktsmuskulaturen
      1 ansiktsnerv
      1 ansiktsnerven
      1 ansiktsområdet
      1 ansiktspiercingar
      2 ansiktsrodnad
      1 ansiktsrörelser
      1 ansiktssjukgymnastik
      1 ansiktssvullnaden
      7 ansiktsuttryck
      1 ansiktsuttrycket
      1 ansiktsvävnad
      1 ansiktuttryck
      1 ansiniso
      1 ansistandard
      1 anskaffade
      3 anslag
      1 anslogs
      1 anslöt
      4 ansluta
      4 anslutande
      1 anslutas
      4 ansluten
      3 ansluter
      1 anslutet
      1 anslutit
      8 anslutna
     25 anslutning
      1 anslutningar
      1 anslutningsmöjligheter
      7 ansluts
      5 ansöka
      6 ansökan
      1 ansöker
      1 ansökningar
      1 ansökningsförfarande
      4 anspänning
      1 anspelar
      6 anspråk
      1 anspråken
      1 anspråkslöshet
      1 anställa
      1 anställas
      7 anställd
     19 anställda
      1 anställde
      1 anställer
      6 anställning
      1 anställs
      1 anställts
      6 anstalt
      1 anstaltref
      1 anständiga
      2 anstränga
      3 ansträngande
      1 ansträngd
      1 ansträngda
      2 anstränger
     20 ansträngning
      1 ansträngningar
      3 ansträngningen
      1 ansträngnings
      4 ansträngningsinkontinens
      2 ansträngs
      1 ansträningsinkontinens
      2 ansvällning
      1 ansvälls
     33 ansvar
      3 ansvara
      1 ansvarade
     24 ansvarar
     16 ansvaret
     15 ansvarig
      9 ansvariga
      1 ansvarsbefriade
      1 ansvarsfull
      1 ansvarslöshet
      1 ansvarslöst
      3 ansvarsområde
      1 ansvarsområdena
      1 ansvarsområdet
     14 anta
      7 antabus
      1 antaga
      5 antagande
      8 antaganden
      1 antagandena
      9 antagandet
      1 antaget
      4 antagit
      4 antagits
     13 antagligen
      1 antagna
      3 antagning
      2 antagonist
      3 antagonisten
      3 antagonister
    218 antal
    182 antalet
      1 antända
      1 antänder
      1 antändningsbar
      1 antänds
     13 antar
      5 antarktis
     47 antas
      1 antecedenter
      1 antecknar
      1 anteckning
      3 anteckningar
      1 anteckningarna
      1 anteckningsbok
      1 antegrad
      1 antenn
      1 antennbärare
      1 antenner
      1 antennerna
      1 anteriort
      1 anterograd
      1 anthelmintikum
      1 anthony
      1 anthophyllum
      2 anthracis
      1 anthrax
      4 anti
      1 antianimaliska
      3 antibakteriell
      8 antibakteriella
      4 antibakteriellt
    183 antibiotika
      1 antibiotikaadministrering
      2 antibiotikaanvändning
      3 antibiotikabehandlade
      1 antibiotikabehandlar
     34 antibiotikabehandling
      2 antibiotikabehandlingar
      1 antibiotikabehandlingen
      1 antibiotikaceftriaxon
      3 antibiotikadosen
      1 antibiotikaförsäljning
      1 antibiotikaförskrivning
      1 antibiotikainjektioner
      1 antibiotikaintag
      1 antibiotikakänsliga
      2 antibiotikakänslighet
      1 antibiotikaklass
      5 antibiotikakur
      2 antibiotikakurer
      1 antibiotikaliknande
      9 antibiotikan
      1 antibiotikaprofylax
     24 antibiotikaresistens
      1 antibiotikaresistensspridning
      1 antibiotikaresistent
      3 antibiotikaresistenta
      1 antibiotikas
      1 antibiotikasalva
      1 antibiotikasorter
      2 antibiotikaterapi
      2 antibiotikatyper
     28 antibiotikum
      1 antibiotikumen
      3 antibiotikumet
      1 antibiotikums
      1 antibiotisk
      2 antibiotiska
      1 antibody
      1 antibodydependent
      1 anticimex
      1 anticipation
      2 antidepressiv
     29 antidepressiva
      1 antidepressivmedel
      3 antidepressivt
      1 antidepressivum
      6 antidiuretiskt
      1 antidopaminerg
      4 antidot
      1 antidotus
      5 antiemetika
      1 antiendomysiumantikroppar
      7 antiepileptika
      1 antiepileptiska
      1 antiepileptiskt
      1 antifosfolipidsyndrom
      1 antifouling
      1 antifrysprodukter
     30 antigen
      1 antigenantikroppkomplex
      2 antigendetektion
      1 antigene
      3 antigenen
     11 antigener
      6 antigenet
      1 antigenetiska
      1 antigenpåvisning
      3 antigenpresenterande
      1 antiglobaliserings
      1 antigraviditetshormon
      1 antihelmintika
      1 antihistamin
      8 antihistaminer
      2 antihistaminpreparat
      1 antihistamintabletter
      1 antihjältar
      1 antihjärna
      1 antihomosexlag
      1 antihomotoxisk
      1 antiigeantikroppen
      1 antiinflamatorika
      8 antiinflammatorisk
     15 antiinflammatoriska
      6 antiinflammatoriskt
      2 antiinflammatory
      1 antiischemiskt
      5 antik
     27 antika
     26 antiken
     15 antikens
      1 antikoagel
      1 antikoagulant
      5 antikoagulantia
      1 antikoagulantiat
      1 antikoagulantium
      1 antikoagulationsmedel
      1 antikoagulatorisk
      2 antikoagulerande
      2 antikolinerga
      2 antikolinergika
      1 antikonvulsivmedicinering
      3 antikropp
     98 antikroppar
      7 antikropparna
      4 antikroppen
      1 antikroppsberoende
      2 antikroppsbildning
      1 antikroppsbildningen
      1 antikroppslösningar
      1 antikroppsproducerande
      2 antikroppsproduktion
      3 antikroppstest
      1 antikroppstitrar
      1 antikroppsutveckling
      1 antikvarisk
      1 antileukotriener
      1 antiloper
      1 antimalariamedel
      1 antimaskmedel
      2 antimikroba
      2 antimikrobiell
      1 antimikrobiella
      1 antimons
      1 antimülleriskt
      1 antimüllerskt
      5 antimykotika
      1 antimykotikaanvänds
      1 antimykotiska
    214 antingen
      1 antinoradrenerg
      1 antinous
      1 antiöstrogena
      6 antioxidant
      4 antioxidanter
      3 antioxiderande
      3 antiparasitära
      1 antiparasitiskt
      1 antipartikel
      1 antipc
      1 antipcnvåer
      1 antipersipranter
      1 antiperspirant
      1 antiperspirantagenser
      1 antiperspirantdeodoranter
      7 antiperspiranter
      1 antiplackbildande
      1 antiprogesteron
      1 antipsykiatri
      4 antipsykiatrirörelsen
      4 antipsykiatriska
      8 antipsykotika
      2 antipsykotikum
      6 antipsykotisk
     12 antipsykotiska
      1 antipyretikum
      1 antiretroviral
      2 antiretrovirala
      2 antireumatiska
      1 antirheumatic
      1 antirökningskampanjen
      3 antirökningskampanjer
      1 antirökningsrörelsen
      1 antirökningsrörelsens
      4 antiseptik
      6 antiseptika
      1 antiseptiken
      3 antiseptikum
      3 antiseptisk
      7 antiseptiska
      7 antiseptiskt
      2 antiserum
     10 antisocial
      1 antisociala
      1 antisocialt
      1 antispasmolytikum
      1 antisvampmedel
      1 antisvettning
      1 antisyfilitiska
      1 antiterrorism
      1 antitnf
      1 antitnfläkemedel
      1 antitransglutaminasantikroppar
      4 antitrombin
      1 antitrombinbrist
      1 ��antitrypsinbrist
      1 antivenom
      4 antiviral
     15 antivirala
      1 antiviralt
      4 antivirusmedel
      1 antivirusmedlet
      1 antivivisektionism
      6 antofyllit
      9 antog
     23 antogs
      6 antoine
      1 antomiska
      4 anton
      3 antonie
      1 antonii
      1 antonitorden
      5 antonius
      5 antoniuseld
     16 antonovsky
      6 antonovskys
     12 antracen
      1 antracenderivat
      1 antracenol
      1 antracenreaktionerna
      1 antracens
      1 antracyklin
      1 anträffats
      2 antrakinon
      1 antrakinonprocessen
      3 antrakos
      1 antrol
      2 antropologen
      1 antropologer
      2 antropologi
      1 antropologin
      1 antropologisk
      1 antroposofi
      1 antroposofin
      3 antroposofisk
      2 antroposofiska
      4 antroposofiskt
      1 antrum
      1 antwerpen
      3 antyda
      2 antydan
      2 antydde
     30 antyder
      1 antydningar
      4 antytt
      1 antytts
      1 anuri
     23 anus
      1 anusarayoga
      1 anusregionen
     19 använd
    255 använda
     11 användande
     32 användandet
     12 användare
     16 användaren
      8 användarens
      1 användarinterfacet
      2 användarna
      1 användarvänligt
    361 användas
     15 användbar
     10 användbara
      2 användbarhet
      2 användbarheten
     17 användbart
     61 använde
    256 använder
    165 användes
    295 användning
      2 användningar
      1 användningarområden
     44 användningen
      3 användningsförbud
      1 användningshistorik
     17 användningsområde
     33 användningsområden
      6 användningsområdet
      1 användningstid
      1 användningstiden
      1 användningstillfälle
   1218 används
     34 använt
    145 använts
      1 anvisning
      3 anvisningar
      1 anvisningarna
      1 anxiolytikum
      1 any
      2 ånyo
     16 aorta
      1 aortaaneurym
     16 aortaaneurysm
      4 aortabågen
      1 aortablodkärl
      1 aortabråck
      3 aortadissektion
      1 aortae
      1 aortakärlet
      5 aortaklaffen
      3 aortan
      1 aortasinus
      1 aortaväggen
      1 aortaväggens
      1 aortit
      1 ap
      3 apa
      1 apan
      1 apas
     14 apati
      2 apatisk
      3 apatiska
      1 apbi
      1 apbibehandling
      1 apd
      1 apdmaskin
      2 apelsin
      2 apelsinhud
      1 aperts
      2 apex
      1 apfonderna
      1 apg
      2 apgar
      1 apgarskalan
      1 apikal
      1 apikalt
      1 apis
      2 aplasia
      1 aplastisk
      3 apné
      6 apnéer
      1 apnéskenor
      1 apnjurar
      1 apodesmos
      1 apodos
      1 apoferritin
      1 apoidae
      1 apokarpa
      1 apoketet
      1 apokrina
      1 apoliva
      1 apollinaire
      3 apollon
      1 apomethyldopa
      1 apomixis
      1 apomorfin
      1 aponno
      1 apoplexi
      9 apoptos
      1 apoptosinducerare
     12 apor
      2 aporna
      1 apostlagärningarna
     30 apotek
     13 apotekare
      3 apotekaren
      1 apotekarens
      1 apotekareverksamhet
      2 apotekarexamen
      1 apotekarlegitimation
      1 apotekarprogrammen
      1 apotekarstudenten
      2 apotekarutbildning
      2 apotekarutbildningen
      2 apotekaryrkena
     12 apoteken
     10 apoteket
      1 apotekets
      1 apoteksassistenter
      1 apoteksbolaget
      1 apoteksgöromål
      1 apotekshandeln
      1 apoteksinstitutionen
      1 apotekskedjan
      2 apoteksmarknaden
      1 apoteksmonopolet
      1 apoteksordningar
      1 apotekspraktik
      1 apotekspraktiken
      1 apoteksprivilegium
      1 apoteksrörelsen
      1 apoteksservicepunkter
      1 apotekstekniker
      1 apotekstillstånd
      1 apoteksvaror
      1 apoteksväsendet
      2 apoteksverksamhet
      1 apoteksverksamheten
      1 apotheke
     13 apparat
     10 apparaten
      1 apparatens
      8 apparater
      1 apparatfelsmodellen
      1 apparatmiljö
      1 apparattyp
      3 apparatur
      1 apparaturen
      1 appeals
      1 äppelcidervinäger
      1 äppelform
      2 äppelformad
      1 appellationsdomstolen
      1 appeller
      4 appendicit
     10 appendix
      2 äpple
      2 äpplen
      1 äpplepäron
      1 appliance
      3 applicera
      1 applicerades
      3 applicerar
     30 appliceras
      1 applicerat
      1 applicerats
      1 applicerbart
      2 applicering
      2 appliceringar
      1 applikation
      1 applikationen
      4 applikationer
      3 applikator
      1 applikatorer
     13 applikatorerna
      1 applikatorernas
      2 applikatorn
      1 apportering
      1 appreteringsprocess
      1 approaches
      1 approximationen
      1 approximativt
     39 apraxi
      1 apraxin
      1 aprd
      1 aprea
      1 aprikos
      1 aprikoser
      1 aprikoskärnor
     22 april
      1 apteksfumar
     11 aptit
      5 aptiten
      2 aptitförlust
      7 aptitlöshet
      1 aptt
      2 aqua
      1 aquam
      2 aquino
      2 aquitaine
      1 aqva
      1 ar
    964 år
      2 �år
      1 år[]
    108 År
  14499 är
     29 Är
      1 ära
      1 arab
      2 araber
      1 araberna
      2 arabicum
      1 arabisk
     11 arabiska
      1 araceae
      1 arachnoidala
      1 arafat
      1 aragonit
      1 araknoidea
      3 åratal
     55 arbeta
     17 arbetade
      1 arbetades
      2 arbetande
    108 arbetar
      1 arbetarbina
      5 arbetare
      1 arbetarfamiljer
      1 arbetarinom
      1 arbetarklasslusken
      5 arbetarna
      1 arbetarrörelsens
      2 arbetarskydd
      1 arbetarskyddsregler
      1 arbetas
      7 arbetat
    123 arbete
     14 arbeten
     51 arbetet
      1 arbetmiljöverket
      4 arbets
      1 arbetsam
      1 arbetsbänkar
      3 arbetsbelastning
      1 arbetsbordet
      1 arbetsdag
      2 arbetsdagar
      2 arbetsdagen
      1 arbetsdefinition
      1 arbetseffekt
      1 arbetsekg
      2 arbetsfält
      1 arbetsförhållanden
      2 arbetsförhållandena
      1 arbetsförlust
      2 arbetsförmåga
      1 arbetsförmågan
      2 arbetsförmedlingen
      1 arbetsgången
     14 arbetsgivare
     11 arbetsgivaren
      4 arbetsgivarens
      1 arbetsgivares
      1 arbetsgivarna
      1 arbetsgivarorganisationerna
      2 arbetsgrupp
      2 arbetsgruppen
      1 arbetsgrupper
      1 arbetsgrupperna
      1 arbetshälsa
      1 arbetshandikapp
      1 arbetshandledning
      1 arbetshjälpmedel
      1 arbetshöjd
      1 arbetsinnehåll
      1 arbetsinsats
      2 arbetskamrater
      1 arbetskapacitet
      4 arbetskläder
      1 arbetsklimat
      2 arbetskostnaden
      1 arbetskraft
      1 arbetskrav
      2 arbetsledare
      2 arbetsliv
     13 arbetslivet
      1 arbetslivets
      1 arbetslivsforskning
      1 arbetslivsinriktad
      1 arbetslivsmuseum
      1 arbetslöhet
      1 arbetslokal
      1 arbetslösa
      6 arbetslöshet
      1 arbetsmängd
      1 arbetsmarknaden
      1 arbetsmaterial
      1 arbetsmetod
     26 arbetsmiljö
      1 arbetsmiljöansvaret
     10 arbetsmiljöarbete
     14 arbetsmiljöarbetet
      1 arbetsmiljöenkäter
      1 arbetsmiljöföreskrifter
      1 arbetsmiljöfrågor
      1 arbetsmiljöhot
      1 arbetsmiljökommissionen
      9 arbetsmiljölagen
      1 arbetsmiljölagstiftningen
     16 arbetsmiljön
      1 arbetsmiljöombud
      1 arbetsmiljöområden
      5 arbetsmiljöpolicy
      1 arbetsmiljöpolicyn
      1 arbetsmiljöproblem
      1 arbetsmiljöproblemet
      1 arbetsmiljörättsliga
      1 arbetsmiljörisker
      1 arbetsmiljöskäl
      8 arbetsmiljöverket
     10 arbetsmiljöverkets
      4 arbetsminne
      3 arbetsminnesträning
      1 arbetsminnesträningsprogrammet
      4 arbetsminnet
      1 arbetsmodeller
      2 arbetsmoment
      1 arbetsnamnet
      1 arbetsoförmåga
      1 arbetsolyckan
      4 arbetsolyckor
      2 arbetsområde
      4 arbetsområden
      1 arbetsområdena
      2 arbetsorganisation
      2 arbetsorganisationen
      1 arbetsorganisationens
      1 arbetsorienterad
      1 arbetspassen
      1 arbetsperioder
      1 arbetsplan
      1 arbetsplanering
     11 arbetsplats
     12 arbetsplatsen
      2 arbetsplatsens
     10 arbetsplatser
      3 arbetsredskap
      1 arbetsrelaterad
      1 arbetsrelaterade
      1 arbetsrelaterat
      1 arbetsresultat
      1 arbetsrock
      1 arbetsroll
      1 arbetssammanhang
      1 arbetssätt
      1 arbetssättet
      2 arbetssituation
      2 arbetssjukdomar
      5 arbetsskada
      2 arbetsskadan
      1 arbetsskadeanmälningar
      4 arbetsskador
      2 arbetsställe
      1 arbetsställning
      6 arbetsställningar
      1 arbetsställningen
      1 arbetsstationer
      1 arbetssuppgifter
      1 arbetssvårigheter
      1 arbetssysslor
     10 arbetstagare
      1 arbetstagaren
      2 arbetstagares
      2 arbetstagarna
      1 arbetstagarnas
      1 arbetstagarorganisationen
      1 arbetstakt
      1 arbetsteknik
      1 arbetstekniskt
      1 arbetstempo
      1 arbetstempot
      9 arbetsterapeut
     13 arbetsterapeuten
      1 arbetsterapeutens
      9 arbetsterapeuter
      1 arbetsterapeuterna
      5 arbetsterapeutiska
      2 arbetsterapeutprogrammet
      1 arbetsterapeututbildningen
     14 arbetsterapi
      1 arbetsterapihuset
      1 arbetsterapin
      7 arbetsterapins
      4 arbetstid
      1 arbetstider
      1 arbetstillfällen
      8 arbetsuppgifter
      2 arbetsuppgifterna
      1 arbetsuppift
      1 arbetsutrustningar
      1 arbetsutrymme
      1 arbiträra
      1 arbovirus
      3 archeus
      1 archie
      1 architecture
      1 archiving
      1 arctica
      1 arcuatus
      1 ard
      2 arden
      1 arderne
      2 ards
      4 are
      2 area
      1 areaktioner
      1 arealer
      1 arean
      2 areata
     75 åren
      2 Åren
      1 arena
      1 arenan
      1 arenaviridae
      3 ärende
      1 ärendehantering
      4 ärenden
      3 ärendet
      1 arenosus
      1 arenreceptorinteragerande
      1 årens
      1 ares
     36 året
      7 Året
      2 aretaeus
      1 årets
      1 arévalos
      1 ärft
     41 ärftlig
     47 ärftliga
      2 Ärftliga
      1 ärftliggenetiskt
     15 ärftlighet
     10 Ärftlighet
      1 ärftligheten
      1 Ärftligheten
      1 ärftlighetens
      1 ärftlighetsfaktorn
      1 ärftlighetsgång
      1 ärftlighetsmönster
      1 ärftligrisken
     17 ärftligt
      2 arg
      2 arga
      2 argentina
      1 argentum
      1 argolis
      1 argon
      1 argos
      1 argt
     16 argument
      4 argumenten
      1 argumentera
      5 argumenterar
      2 argumenterat
      2 argumenterats
      2 argumentet
      1 argyll
      7 århundrade
      6 århundraden
      3 århundradena
      6 århundradet
      1 Århus
      1 aria
      1 arianska
      2 aricept
     15 årig
      2 åriga
      3 årige
      1 arillus
      3 åringar
      1 åringars
     18 aripiprazol
      2 aripiprazole
      4 ariska
      1 aristokrater
      1 aristokratiskt
      2 aristolochia
      9 aristoteles
      1 arizonicus
      1 arjeplogssjukan
      1 arjohuntleigh
      3 ark
      1 arkansas
      1 ärkebiskop
      4 arkebusering
      1 ärkedum
      1 arkéer
      1 arkeologen
      2 arkeologer
      1 arkeologi
      2 arkeologisk
      3 arkeologiska
      2 arkeo�logiska
      1 arketyper
      1 arkitekter
      1 arkitektur
      1 arkitekturen
      1 arkitekturer
      1 arkiv
      1 arkiveras
      4 arktis
      1 arktiska
      1 arkuatuskärnan
      5 årlig
     10 årliga
     43 årligen
      4 Årligen
     23 arm
      1 armani
     29 armar
      1 ärmar
     12 armarna
      2 armauer
      1 armbågar
      6 armbågen
      4 armbågens
      1 armbågsled
      1 armbågsleder
      1 armbågslederna
      1 armbågsledsartros
      3 armbågsledsdysplasi
      2 armé
      2 arméer
      1 arméerna
      1 arméknivar
     17 armen
      7 armén
      1 armeniska
      2 arméns
      1 armenus
      1 armera
      1 armeras
      2 armering
      5 armhålan
      1 armhåle
      8 armhålor
      5 armhålorna
      2 armillaria
      1 armkläde
      1 armlängd
      1 armleden
      1 armmageskinka
      1 armmovement
      1 armproteser
      1 armrörelser
      1 armstyrka
      1 armveck
      1 armvecken
      2 armvecket
      1 arne
      2 arnica
      1 arnicadrogen
      1 arnicadrogerna
      3 arnicae
      1 arnikor
      1 arnims
      2 arnold
      1 arnoldchiaris
      2 äro
      2 ärofullt
      1 arom
      1 aromalampor
      1 aromämnen
      3 aromatas
      1 aromatasbrist
      1 aromatashämmande
      2 aromatashämmare
      1 aromaterapi
      1 aromaticitet
      1 aromatisering
      8 aromatisk
      5 aromatiska
      7 aromatiskt
      2 aromer
      2 arousal
     20 ärr
      2 ärrad
      3 arrangemang
      5 arrangera
      1 arrangerade
      1 arrangerandet
      1 arrangerat
      8 ärrbildning
      3 ärrbildningar
      1 ärrbildningen
      1 ärrbråck
      2 ärren
      1 Ärren
      1 arrestlokal
      1 ärret
      1 arrhenius
      6 ärrvävnad
      1 ars
    154 års
     24 årsåldern
      3 �årsåldern
      1 årsarbetstid
      1 årsbasis
      1 årsbehovet
      1 arsea
      1 arsenal
      2 arsenicum
      1 arsenider
     26 arsenik
      2 arseniken
      1 arsenikens
      1 arsenikföreningar
      1 arsenikföreningen
      2 arsenikförgiftning
      1 arsenikinnehållande
      1 arsenikjärn
      2 arsenikkis
      1 arsenikon
      1 arsenikorganiskt
      1 arsenikpentoxid
      1 arseniksulfid
      1 arseniktriklorid
      6 arseniktrioxid
      9 arsfenamin
      1 arsfenaminsalvarsan
      1 årsgrupperna
      1 arsinoe
      2 årsjubileum
      1 årsöverlevnaden
      2 årsperiod
      1 årsredovisningen
      1 årsringar
      2 årsskiftet
      3 årsskott
      4 årstid
      3 årstiden
      1 årstider
      1 årstiderna
      1 årstidsbunden
      1 årstidsbundet
      1 årstidsvariationer
      2 Årsunda
     93 art
      1 ärt
      3 ärta
      1 ärtajordnötsoja
      1 årtal
      1 artantal
     14 artär
      1 artärblodets
      2 artärbråck
      1 artäremboli
      4 artären
      1 artärens
     27 artärer
      5 artärerna
      2 artärernas
      1 artärgren
      1 artäriell
      1 artärinflammation
      1 artäriska
      1 artärsidan
      1 artärskada
      1 artärspasm
      1 artärt
      1 artärvolymer
      1 artefakt
      2 artefakter
     91 arten
      7 artens
      1 artepitet
      3 artepitetet
    177 arter
      1 ärter
      4 arteria
     11 arteriell
      3 arteriella
      3 arteriellt
      1 arteriografi
      1 arteriol
      1 arteriolens
      3 arterioler
      1 arteriolerna
      1 arteriolernas
      6 arterioskleros
      1 arteriöst
      1 arteriosus
      2 arteriovenös
      1 arteriovenösa
      1 arterit
     33 arterna
      1 arternas
      2 arteroskleros
      1 arters
      1 artfränder
      1 artgränser
      1 artheroskleros
      1 arthron
      6 arthur
      1 artiell
      2 artificiell
      3 artificiella
      6 artificiellt
     33 artikel
     23 artikeln
     15 artiklar
      3 artiklarna
      3 artikulation
      2 artikulationen
      1 artikulationsapraxi
      1 artikulationsrörelser
      1 artikulera
      1 artikulerat
      2 artilleri
      2 årtionde
      6 årtionden
      2 årtiondena
      3 årtiondet
      1 årtiondets
      1 artist
      2 artisten
      3 artister
      1 artistnamn
      2 artnamnet
      2 arton
      1 artonårsåldern
      2 artonde
      1 ärtor
      1 artoskop
      1 artoskopet
      4 artralgi
      1 art�ria
      1 art�riae
      2 artrikt
     27 artrit
      2 artriten
      5 artriter
      1 artritsjukdomar
      2 artrodes
      2 artropati
      1 artropatier
      1 artropatierna
     13 artros
      2 artrosen
      1 artroskopi
      1 artrosledförslitning
      1 artrossjukdomarna
      1 arts
      1 artspecifika
      2 artur
      3 årtusenden
      7 ärtväxter
      1 årundradet
     20 arv
      3 ärva
      3 ärvas
      1 ärvda
      1 ärvde
      4 ärver
      1 arvet
      2 arvid
      1 arvo
      1 arvprinsen
     11 ärvs
      6 arvsanlag
      2 arvsanlagen
      1 arvsberoende
      8 arvsmassa
      9 arvsmassan
      1 arvsmassans
      1 arvsrätt
      4 ärvt
      1 arvtagaren
      1 ärvts
      1 arybrosk
      1 aryl
      1 arytenoidea
      7 arytmi
      1 arytmibenägenhet
     10 arytmier
      1 arytmierna
      1 arytmin
      1 ärztlichen
     12 as
      1 ås
      1 Äs
      2 asa
      2 Åsa
      1 asacol
      3 asainducerad
      1 åsamka
      1 åsamkar
      1 åsamkas
      1 äsan
      3 asana
      2 asanas
      2 åsar
      2 asas
      1 asasbindningar
      6 asat
      2 asatalatkvot
      2 asätare
      1 Åsberg
     70 asbest
      2 asbestanvändning
      7 asbestcement
      1 asbestcementledningar
      3 asbestcementplattor
      2 asbestcementrör
      1 asbestcementskivor
      7 asbestexponering
      1 asbestfiber
     15 asbestfibrer
      1 asbestfibrerna
      1 asbestfibrernas
      1 asbestfibrers
      1 asbestfri
      1 asbestfria
      5 asbesthaltiga
      3 asbesthaltigt
      1 asbestisolering
      3 asbestmaterial
      1 asbestmaterialen
      6 asbestmineral
      1 asbestmineralet
      3 asbestorsakade
     16 asbestos
      1 asbestprevention
      1 asbestproducerande
      1 asbestrelaterad
      2 asbestrelaterade
      2 asbestsanering
      2 ascaris
      1 aschheim
     19 ascites
      1 ascitesvätskan
      1 ascl
      1 ascosporer
      5 asd
      5 aseptik
      1 aseptiken
      3 aseptikens
      6 aseptisk
      2 aseptiskt
      1 åser
      1 asexualitet
      6 asexuell
      1 asexuella
      7 asexuellt
      1 asfalt
      1 asfalten
      1 asfaltlim
      1 asfaltsrester
      1 asfäriska
      1 asfyktiska
      1 asfyxi
      1 ashermans
      2 ashtanga
      1 ashtangas
      1 ashtangayoga
      1 ashvinerna
      1 asia
      1 asiaten
      2 asiater
      3 asiatisk
      7 asiatiska
      2 asiatiskt
      1 åsidosätta
      1 åsidosättande
     65 asien
      4 åsikt
      1 åsikten
      9 åsikter
      2 åsikterna
      1 asimov
      2 ask
      1 aska
      2 åska
      1 åskådare
      4 åskådliggör
      1 åskådliggöra
      1 åskådning
      1 askar
      1 askarna
      1 asketer
      1 asketiska
      1 asketism
      2 askfat
      1 åskguden
      1 askitesvätska
      2 asklepeia
      3 asklepiades
     13 asklepios
      1 asklepiosstaven
      1 asklut
      3 askorbinsyra
      1 asks
      1 askträd
      1 åskvigg
      1 Åsling
      1 asmatstammarna
      1 Åsmund
      1 åsna
      1 åsninna
      2 åsnor
      2 aso
      3 asociala
      1 aspartat
      1 aspartataminotransferas
      8 aspekt
      3 aspekten
     25 aspekter
      3 aspekterna
      2 asperger
      1 aspergerliknande
     14 aspergers
      1 aspergillom
      4 aspergillos
      2 aspergillus
      1 aspergillussporer
      1 aspergillussvampen
      1 aspermi
      1 asphyxia
      1 aspidogastrea
      6 aspiration
      1 aspirationbrus
      1 aspirationen
      1 aspirationer
      7 aspirationspneumoni
      1 aspirationspneumonit
      1 aspirera
      3 aspirerade
      2 aspirerar
      1 aspirerat
      3 aspirin
      1 asplund
      1 asrashexahydrometoximetylah[]bensofuro[aef]
      3 assay
      1 assemblerkod
      1 assemblerspråk
      2 assembly
      1 assertive
      2 assesment
      1 assimilationer
      1 assimileras
      1 assimilerats
      1 assimilering
      2 assistance
      2 assistans
      1 assistanshundarna
      1 assistanshunden
      1 assistant
      2 assisted
      4 assistent
      2 assistenter
      2 assistera
      6 assisterad
      1 assisterade
      2 assisterar
      2 assisterat
      3 associated
     23 association
      3 associationer
      1 associationerna
      2 associations
      4 associationsbesvär
      1 associationskärnor
      1 associationsstudier
      4 associera
      5 associerad
     24 associerade
      1 associerades
      3 associerar
     20 associeras
     14 associerat
      4 associerats
      1 asss
      1 assumption
      1 assyrien
      1 assyrier
      2 assyriska
      3 ast
      3 åstadkom
     20 åstadkomma
      6 åstadkommas
      7 åstadkommer
      3 åstadkommes
      2 åstadkoms
      1 astaxantin
      5 asteni
      1 asterisk
      1 asterixis
      1 asthanga
      1 asthi
      2 asthma
      3 astigmatism
     68 astma
      1 astmaanfall
      1 astmaattack
      1 astmaattacker
      2 astmabehandling
      1 astmabesvär
      1 astmaexacerbationer
      2 astmaförsämringar
      2 astmakontroll
      1 astmaläkemedel
      1 astmaliknande
      1 astmamediciner
      1 astman
      2 astmasymtom
      1 astmatest
      6 astmatiker
      1 astmatiska
      1 astmatiskt
      1 astomi
      3 astra
      1 astral
      2 astralkropp
      1 åstränder
      1 astreptokocker
      2 astrid
      1 astrocytens
      4 astrocyter
      4 astrocyterna
      1 astrocytom
      2 astrocytutskott
      1 astrocytutskotten
      1 astrofysik
      2 astronauter
      2 astronomi
      2 astronomin
      1 astronomiska
      1 åsyfta
      2 åsyftade
      8 åsyftar
      4 åsyftas
      2 asyler
      1 asylinrättningarna
      3 asymmetrisk
      7 asymptomatisk
      2 asymptomatiska
      1 asymptotiskt
      9 asymtomatisk
      4 asymtomatiska
      3 asymtomatiskt
      1 asystemet
      2 asystoli
      5 at
    187 åt
      1 Ät
     92 äta
      2 åtagande
      2 åtaganden
      1 åtagit
      1 ataktisk
      4 åtal
      3 åtalad
      2 åtalade
      3 åtalades
      1 atanatologi
      6 ätande
      1 åtanke
     16 ätas
      7 ataxi
      1 ataxier
      1 ataxisjukdomar
      1 ataxisjukdomen
      5 ätbara
      1 ätbegär
      1 ätbeteendet
      1 åtbörder
      4 atc
      2 atcantenn
      1 atcbesked
      1 atcfel
      1 atckod
      1 atckoden
      3 atcsystemet
      1 åtdraget
      1 åtehämtar
      1 ateism
      1 ateister
      2 atelektas
      2 atelektaser
      1 ateles
      3 aten
      1 äten
     24 åter
      2 Åter
     91 äter
      2 Äter
      2 återabsorberas
      1 återandningsteknik
      1 återanpassa
      1 återanslutas
      1 återanvända
      5 återanvändas
      1 återanvändningsbar
      3 återanvändningsbara
      1 Återanvändningsbara
      2 återanvänds
      1 återberättar
      1 återberättats
      3 återbesök
      1 Återbesöken
      2 återbilda
      6 återbildas
      4 återbildning
      1 återbyggnadsprocessen
      1 återdraperas
      7 återfå
     16 återfall
      1 Återfall
      1 återfallen
      1 återfaller
      1 återfallsfeber
      1 återfallsförbrytare
      1 återfallsfritt
      1 återfallsprevention
      1 återfallsrisken
      2 återfanns
      4 återfår
      2 återfås
      1 återfått
      1 återfinna
      7 återfinnas
      1 återfinner
     53 återfinns
      1 återfjädringstryck
      3 återflöde
      4 återflödet
      2 återfödas
      3 återfödelse
      2 återfödelsen
      1 återfödelsens
      1 återfödelser
      3 återföds
      1 återföll
      1 återför
      3 återföra
      2 återföras
      1 återförenas
      2 återförs
      2 återförsäljare
      1 återfukta
      1 återfunnen
      6 återfunnits
     12 återgå
      1 återgången
     11 återgår
      1 återgått
      4 återge
      1 återger
      1 återgetts
      1 återgick
      1 återgivas
      1 återgivits
      1 återgivning
      1 återgivningar
      1 återhållsamhet
      4 återhämta
      7 återhämtar
      3 återhämtat
     13 återhämtning
      4 Återhämtning
      3 återhämtningen
      1 återhämtningsfas
      1 återhämtningsgrupper
      1 Återhämtningsprojektet
      1 återhämtningstiden
      1 Återhämtningstiden
     15 återigen
      1 Återigen
      1 återinfektion
      1 återinfektioner
      2 återinföra
      1 återinförandet
      1 återinförts
      1 återinsjuknande
      1 återintroduceras
      1 återinvesteras
      2 återkallas
      4 återkom
     11 återkomma
     51 återkommande
      4 Återkommande
     21 återkommer
      2 återkommit
      3 återkomsten
      1 återkoppla
      1 återkoppling
      1 återkopplingstakykardier
      1 återlämnas
      2 aterom
      1 återomvandlas
      9 ateroskleros
      1 aterosklerotiskt
      1 återprojektion
      1 återrapportering
      1 återsända
      7 återskapa
      2 återskapande
      1 återspegla
      7 återspeglar
      1 återspeglas
      3 återstående
     18 återställa
      6 återställd
      3 återställer
      8 återställs
      3 återstår
      1 återstoden
      1 återsuget
      1 återta
      1 återtagande
      1 återtagandet
      2 återuppbyggnad
      1 återuppfödningssyndrom
      2 återupplevande
      1 återupplevandesymtom
      1 återupplivningsresultat
      1 återupprätta
      1 återupprepade
      1 återuppstå
      1 återuppståndelse
      1 återuppstått
      2 återuppstod
      1 återupptag
      4 återupptaget
      2 återupptas
      3 återupptogs
      1 återuppväcka
      1 återuppväckt
      1 återuppväcktes
      1 återuppvärms
      1 återväcktes
      1 Återvänd
      6 återvända
      1 återvändande
      4 återvände
      6 återvänder
      1 återvanns
      3 återvänt
      1 återväxten
      1 återverkningar
      1 återvinnas
      1 återvinningsbar
      1 återvinningsbara
      1 återvinningsbart
      1 återvinningscentral
      1 återvinns
      1 återvunnen
      5 åtföljande
      3 åtföljas
      1 åtföljd
      1 åtföljda
      1 åtföljer
      4 åtföljs
      1 åtföljt
      2 åtgår
     15 åtgärd
     14 åtgärda
      1 åtgärdades
     12 åtgärdas
      5 åtgärden
    108 åtgärder
     12 Åtgärder
      8 åtgärderna
      1 åtgärdsarbete
      1 åtgärdsförslag
      1 åtgärdsmekanism
      1 Åtgärdsplanen
      1 atharvaveda
      1 Åthävaden
      1 athena
      1 athenaios
      1 athens
      1 athere
     14 ätit
      1 ätits
      7 atkins
      1 atkinsdiet
     13 atkinsdieten
      3 atkinsmetoden
      2 åtkomligt
      4 åtkomst
      1 atl
      2 atläkare
      1 atlantica
      1 atlantiska
      1 atlas
      1 atlaser
      3 ätlig
      8 ätliga
      1 Ätlighet
      2 atm
      1 atma
      8 atman
      1 atmanbrahman
      1 atmans
     56 åtminstone
      3 Åtminstone
      8 atmosfären
      1 atmosfäriskt
      1 atmosfärluft
      2 atmosfärstryck
      1 atnalet
      1 åtnjuter
      1 atÖ
      1 atom
      1 atombombsdetonation
      1 atomen
      4 atomer
      1 atomernas
      1 atomkärnor
      4 atomnummer
      2 atomnumret
      2 atomo
      1 atomoxetin
      1 atomtidsskalan
      1 atomubåtar
      5 atomur
      1 atomuret
      3 atopi
      2 atopisk
      3 atopiska
      3 atopiskt
      1 atorvastatin
      1 atoxyl
     11 atp
      2 åtrå
      1 atralgi
      1 atransferrinemi
      1 åtråvärt
      4 atrazin
      1 atreceptorn
      1 atresi
      1 atretiska
      1 atria
      1 atributen
      2 atrioventrikulära
      8 atrofi
      1 atrofier
      3 atrofisk
      2 atropa
      1 atropatanus
      1 atrophia
      7 atropin
      1 atropos
      3 åts
      9 äts
      3 åtsittande
      3 åtskilda
      8 åtskilliga
      1 Åtskilliga
      2 åtskilligt
      3 åtskillnad
      1 åtskilt
      1 åtsnörd
      6 ätstörning
      2 Ätstörning
     16 ätstörningar
      3 Ätstörningar
      2 ätstörningarna
      1 ätstörningen
      1 ätstörningsdiagnoserna
      1 ätstörningspatienter
  15358 att
     58 åtta
      1 Åtta
      2 åttaårig
      4 attachment
      3 attacin
     11 attack
     14 attacken
     20 attacker
      3 attackera
      3 attackerade
      4 attackerar
     12 attackerna
      3 attackvis
      1 attentat
      5 attention
      1 attenuated
      1 attenuerad
      2 attenuerade
      1 attenueras
      1 attgöralistor
      1 ättika
      1 ättiksinläggning
     16 ättiksyra
      1 ättiksyraanhydrid
      1 ättiksyrans
      1 attila
      3 attityd
      6 attityder
      1 attjänst
      1 ättling
      1 åttlingar
      5 åttonde
      1 åttondelar
      1 åttondels
      1 attract
      1 attraherad
      1 attraherande
      5 attraherar
      2 attraheras
      1 attraherat
      2 attraktion
      2 attraktionen
      1 attraktiv
      4 attraktiva
      1 attraktivitet
      1 attraktiviteten
      4 attraktivt
      1 attrapper
      1 attribueras
      3 attribut
      1 attsocialstyrelsen
      1 atutbildning
      1 ätvanor
      6 atypisk
     18 atypiska
      2 atypiskt
      1 aubrey
      2 audio
      1 audiofrekvenser
      3 audiogram
      2 audiologi
      1 audiologin
      1 audionom
      1 audionomer
      2 audiosignal
      1 audit
      1 auditiv
      6 auditiva
      1 auditivt
      1 audrey
      1 auer
      1 auerstav
      1 auf
      3 auffenberg
      1 auffenbergsexpeditionen
      1 auffenbergsexpeditionens
      3 aufguss
      1 augit
      1 augmented
      5 august
      1 augusta
      1 augustenbad
     20 augusti
      1 augustioktober
      1 augusto
      1 augustus
      1 auktionshusen
      4 auktorisation
      1 auktoriserad
      4 auktoriserade
      1 auktoriserat
      1 auktoritär
      3 auktoritet
      1 aum
      1 aumsekten
      3 aura
      1 auraminrhodaminfärgning
      4 auran
      1 aureolus
     25 aureus
      1 auriculoterapeutiska
      3 auriculoterapi
      3 auror
      5 auschwitz
      3 auskultation
      1 auskultera
      1 austrailien
      1 austral
      2 australia
      4 australian
     46 australien
      3 australiens
      2 australiensisk
      3 australiensiska
      1 australisk
      1 autentisk
      1 authorisation
      1 authority
     86 autism
      1 autismautismliknande
      1 autismbegreppet
      2 autismen
      1 autismens
      3 autismliknande
      1 autismspektra
      1 autismspektrumbegreppet
      3 autismspektrumet
     18 autismspektrumstörning
      3 autismspektrumstörningar
     16 autismspektrumtillstånd
      1 autistischen
      8 autistiska
      8 autistiskt
      1 autoamputation
      1 autoanamnes
      9 autoantikroppar
      1 autofagi
      1 autofagocytos
      1 autofire
     23 autoimmun
     34 autoimmuna
      2 autoimmune
     17 autoimmunitet
      2 autoimmuniteten
      2 autoimmunitetens
      2 autoimmunt
      3 autoinjektor
      3 autoinjektorn
      2 autoklav
      2 autoklaven
      2 autoklaver
      2 autoklavering
      1 autoklavprocessen
      5 autokommunikation
      1 autokorrelationsfunktion
      1 autokrin
      3 autolog
      2 automatic
      3 automatik
      1 automatisera
      1 automatiserad
      3 automatiserade
      1 automatiseras
      1 automatisering
     10 automatisk
      3 automatiska
     20 automatiskt
      6 autonom
     12 autonoma
      2 autonomi
      1 autonomin
      1 autonomt
      1 autopilot
      2 autoregressiv
      1 autos
      1 autosom
      6 autosomalt
      2 autosuggestion
      1 autstraliensiska
      1 autumn
      2 autumnale
      1 auxiner
  16231 av
      2 äv
      2 ava
      3 avägd
      2 availability
      1 avaktivera
     18 avancerad
     19 avancerade
      1 avancerat
      1 avantasia
      1 avantgardistisk
      1 avantgardistiska
      1 avarter
      5 avbilda
      1 avbildade
      1 avbildades
      1 avbildande
      1 avbildandet
      4 avbildar
      6 avbildas
      1 avbildats
      8 avbildning
      1 avbildningarna
      1 avbildningskvalité
      1 avbildningsmetoder
      1 avbildningsteknik
      1 avbildningstekniker
      1 avblir
     14 avblock
      1 avböjda
      1 avböjes
      1 avböjt
      1 avbröts
     12 avbrott
      1 avbrottssjuka
      5 avbruten
      1 avbrutet
      2 avbrutits
      1 avbrutna
      1 avbryt
     10 avbryta
      5 avbrytande
      1 avbrytandet
      6 avbrytas
      5 avbryter
      6 avbryts
     10 avdelning
      8 avdelningar
      1 avdelningarna
      3 avdelningen
      5 avdöda
      1 avdödade
      1 avdödande
      1 avdödar
      1 avdödas
      1 avdödats
      2 avdödning
      2 avdomning
      1 avdragbar
      1 avdunsta
      3 avdunstar
      1 avdunstat
      2 avdunstning
      1 avdunstningen
      1 avdustningen
      6 avel
      1 avelsprogram
   2263 även
    340 Även
      1 avenin
      1 Ävenså
      1 äventyr
      1 äventyrar
      2 avenue
      3 aversion
      1 aversionsterapi
      1 aversiva
      1 avery
      1 avf
      6 avfall
      1 avfallen
      6 avfallet
      1 avfallsämnen
      1 avfallshantering
      1 avfallshink
      1 avfallsmängder
      1 avfallsprodukt
      3 avfallsprodukten
      5 avfallsprodukter
      1 avfärd
      1 avfärdar
      1 avfärdat
      1 avfärgats
      1 avfettande
      1 avfettningssammanhang
      2 avfistel
      1 avflackade
      1 avflackas
      2 avflöde
      1 avflödeshinder
      3 avförande
      1 avförda
     54 avföring
      1 avföringarna
     29 avföringen
      2 avföringens
      1 avföringsfläck
      1 avföringsfläcken
      2 avföringsinkontinens
      1 avföringsinkontinensanalinkontinens
      1 avföringslevande
      2 avföringsmedel
      2 avföringsprov
      1 avföringsprover
      1 avfuktning
      1 avfyra
      1 avfyras
      1 avgå
      1 avgång
      1 avgångsförhör
      5 avgår
      2 avgaser
      1 avgaserna
      1 avgasrening
      2 avgav
     12 avge
     16 avger
      6 avges
      2 avgift
      3 avgifta
      1 avgiftade
      1 avgiftar
      1 avgifter
      3 avgiftning
      1 avgiftsfinansierad
      1 avgiftsfri
      2 avgiftsfria
      1 avgivit
      2 avgjuten
      1 avgjutning
      1 avglottis
     14 avgör
     35 avgöra
     33 avgörande
      1 avgörandet
      4 avgöras
     10 avgörs
      1 avgränsa
      3 avgränsad
      1 avgränsade
      1 avgränsar
      1 avgränsas
      2 avgränsat
      4 avgränsning
      2 avgränsningarna
      1 avgudar
      1 avhållas
      2 avhåller
     14 avhållsamhet
      1 avhämning
      1 avhandlar
      1 avhandlas
     14 avhandling
      4 avhandlingar
      4 avhandlingen
      1 avhängig
      1 avhängiga
      1 avhärda
      1 avhela
      1 avhinfluenzae
      3 avhjälpa
      1 avhjälpande
      2 avhjälpas
      3 avhjälps
      1 avhugget
      1 avhuggning
      1 aviär
      3 avicenna
      1 avicennas
      1 avidin
      1 avigan
      1 avignon
      1 åvilara
      2 avirus
      2 avitamin
      1 avitaminbrist
      3 avium
      1 avkall
      1 avklarad
      1 avklarar
      1 avklinga
      1 avklingande
      2 avklingar
      1 avklipper
      1 avklippta
      1 avknäppbara
      2 avknoppas
      3 avknoppning
      1 avknuta
      9 avknutan
      4 avkoda
      1 avkodning
      1 avkodningen
      1 avkodningsprocessen
      3 avkok
      1 avkomling
      4 avkomlingar
      1 avkomlingarna
     10 avkomma
      7 avkomman
      6 avkommor
      1 avkoppling
      1 avkopplingsfri
      1 avkriminaliserades
      1 avkriminaliserat
      2 avkriminaliserats
      2 avkriminalisering
      1 avkriminaliseringen
      1 avkroka
      1 avkylda
      2 avkylning
      1 avl
      1 avla
      2 avlade
      1 avlades
      1 avlagd
      3 avlägga
      2 avlagringar
      2 avlägsen
      1 avlägset
     48 avlägsna
      2 avlägsnad
      3 avlägsnade
      2 avlägsnades
     10 avlägsnande
      3 avlägsnandet
     10 avlägsnar
     39 avlägsnas
      1 avlägsnat
      6 avlägsnats
      7 avlagt
      1 avlagts
      2 avlång
      1 avlånga
      1 avlänkas
      2 avlänkning
      2 avlänkningen
      1 avlänkningsplattorna
      1 avlar
      8 avläsa
      3 avläsas
      4 avläser
      2 avläsning
      1 avläsningar
      1 avläsningarna
      1 avläst
      3 avlasta
      1 avlastande
      2 avlastas
      1 avläste
      5 avlastning
      2 avlat
      1 avlaten
      1 avlats
     23 avled
      1 avleda
      1 avledare
      1 avledda
      3 avledning
      7 avledningar
      7 avledningarna
      3 avlida
      3 avliden
     14 avlider
      1 avlidet
     10 avlidit
      5 avlidna
      2 avlidne
      3 avliva
      2 avlivas
      2 avlivning
      2 avlönad
      3 avlopp
      1 avloppet
      1 avloppsledningar
      1 avloppsreningsverk
      1 avloppsreningsverket
      2 avloppssystem
      1 avloppsvatten
      6 avloppsvattnet
      1 avlossade
      1 avlossningstillfället
      2 avlövningsmedel
      1 avlunginfiltratlunginflammation
      2 avlusning
      1 avlyssningen
      2 avmagring
      2 avmaskas
      1 avmaskning
      1 avnaprapater
      1 avnjutas
      1 avokado
      1 avokadoolja
      1 avolition
      3 avpassad
      1 avpu
      2 avr
      2 avråda
      2 avrådde
      5 avråder
      4 avråds
      1 avrätta
      1 avrättad
      2 avrättade
      1 avrättas
      4 avrättning
      5 avrättningar
      2 avrättningen
      1 avrättningsgas
      9 avrättningsmetod
      1 avrättningsmetoden
      1 avrättningsprocedurer
      2 avregistrerades
      1 avregistrerat
      2 avreglerades
      1 avregleras
      1 avregleringen
      1 avrinningsområden
      1 avrivningar
      1 avrt
      1 avrundat
      4 avsåg
      2 avsäger
      1 avsågs
      1 avsagt
     42 avsaknad
      8 avsaknaden
      1 avsatt
      1 avsätta
      2 avsatte
      1 avsätter
      1 avsätts
     10 avse
     28 avsedd
     29 avsedda
     31 avseende
      8 avseenden
      1 avseendet
     46 avser
      1 avsersion
     37 avses
     12 avsett
      6 avsevärd
      3 avsevärda
     24 avsevärt
      1 avsides
     10 avsikt
      4 avsikten
      2 avsikter
      1 avsikterna
      2 avsiktlig
      1 avsiktliga
      7 avsiktligt
     11 avskaffades
      2 avskaffandet
      2 avskaffas
      3 avskaffat
      3 avskärmad
      1 avskärmat
      2 avskärmning
      1 avskedsbrev
      2 avskild
      3 avskilda
      1 avskildhet
      2 avskilja
      1 avskiljning
      6 avskiljs
      1 avskilt
      2 avskräcka
      3 avskräckande
      1 avskräcker
      1 avskrevs
      1 avskriva
      1 avskuren
      1 avskurna
      2 avsky
      1 avskydda
      1 avskyvärt
      1 avslå
      1 avslag
      1 avslagna
      1 avslappnade
      1 avslappnande
      1 avslappnat
      4 avslappning
      1 avslappningsövningar
      6 avslöja
      1 avslöjad
      1 avslöjanden
      1 avslöjandet
      6 avslöjar
      3 avslöjas
      1 avslöjat
      6 avsluta
      8 avslutad
      3 avslutade
      2 avslutades
      4 avslutande
      2 avslutar
     24 avslutas
      9 avslutat
      8 avslutats
      1 avslutningen
      2 avsmalnande
      4 avsnitt
      4 avsnittet
      3 avsöndrar
      2 avsöndras
      1 avsöndringen
      1 avsötning
      6 avspänning
      1 avspänningen
      1 avspänningsmetod
      1 avspänningsträning
      2 avspänt
      2 avspärrning
      1 avspegla
      6 avspeglar
      2 avspjälkningen
     17 avstå
     34 avstånd
     14 avståndet
      1 avståndsmarkeringar
      2 avståndssynskärpan
      2 avståndstagande
      1 avstängd
      3 avstängning
      2 avstanna
      2 avstannar
      2 avstannat
      9 avstår
      1 avstavning
      1 avstigmatisera
      2 avstötning
      1 avstötningsreaktion
      2 avstötningsreaktioner
      1 avstötningsrisk
      1 avstressande
      1 avstyra
      1 avsvällande
      1 avsvällning
      1 avsvalnat
      2 avsvalning
      1 avsvära
      1 avsvärande
      1 avsvärtad
      1 avsvärtning
      6 avta
      1 avtäckning
      3 avtagande
      1 avtagbara
      2 avtagit
     10 avtal
      1 avtala
      3 avtalet
      1 avtalsfråga
      1 avtändningen
     13 avtar
      1 avteckna
      1 avtecknade
      2 avtog
      2 avträdet
      1 avtrappning
      4 avtrubbad
      1 avtrubbade
      1 avtrubbning
      1 avtryck
      1 avund
      3 avvägning
      1 avvägningar
      2 avvakta
      1 avvaktan
      1 avvaktande
      3 avvänjning
      1 avvärja
      1 avvärjar
      1 avvärjningsrörelser
      1 avvattna
      1 avvattnade
      1 avvattnas
      1 avvattning
      2 avvecklades
      2 avvecklats
      3 avveckling
      2 avvecklingen
      1 avvek
      2 avverkning
      1 avvika
     36 avvikande
      2 avvikare
     22 avvikelse
      5 avvikelsen
      1 avvikelsens
     26 avvikelser
      1 avvikelserna
      6 avviker
      1 avvisad
      1 avvisade
      1 avvisades
      1 avvisande
      5 avvisar
      2 avvisas
      2 avvisats
      1 avyttrades
      1 award
      2 awareness
      1 away
      1 ax
      5 axel
      5 axelband
      3 axelbanden
      2 axelbandslös
      1 axellångt
      7 axeln
      1 axelns
      2 axelryckning
      1 axelsons
      2 axelsson
      1 axen
      1 axial
      1 axialt
      1 axiella
      1 axiomatisk
      2 axis
      1 axl
     10 axlar
      5 axlarna
      5 axolotl
      1 axolotlen
      6 axon
      1 axonal
      6 axonen
      1 axonens
      3 axoner
      1 axonerna
     13 axonet
      1 axonets
      1 axonterminalen
      1 axoplasmatiskt
      1 ayscough
      1 ayu
     15 ayurveda
      1 ayurvedapreparat
      1 ayurvedaprodukter
      1 ayurvedautbildad
     11 ayurvedisk
      5 ayurvediska
      2 ayus
      1 azatioprin
      1 azedarach
      2 azeotrop
      1 azithromycin
      2 azitromax
      5 azitromycin
      1 azobensen
      1 azofärgämne
      2 azofärgämnen
      1 azoföreningar
      2 azoospermi
      1 azotemi
      5 aztekerna
      3 aztekiska
    117 b
      1 bä
      1 baal
      1 bab
      1 babbage
      1 babianer
      1 babianerna
      1 babianhannen
      1 babraham
      9 baby
      4 babyboom
      1 babyboomgeneration
      1 babycenter
      2 babylonien
      1 babylonier
      1 babylonierna
      1 babyloniska
      1 babyolja
      3 babypuder
      1 babyrytmik
      2 babysim
      1 babyspråk
      3 baccata
      1 bachelor
      1 bachylobum
      1 bacill
      2 baciller
      1 bacillhärdar
      8 bacillus
      1 back
      1 backa
      3 backar
      1 bäckar
      1 backarna
      1 backe
      5 backen
      8 bäcken
      2 bäckenbotten
      3 bäckenbottenmuskulaturen
      2 bäckenbottenövningar
      1 bäckenbottens
      2 bäckenbottenträning
      1 bäckenbottnen
      1 bäckenbottnens
     12 bäckenet
      5 bäckenets
      1 bäckenfogen
      2 bäckenförträngning
      1 bäckenfrakturer
      2 bäckenhåla
      1 bäckenhålan
      1 bäckeningången
      1 bäckenkanalen
      1 bäckenklyvning
      1 bäckenlederna
      2 bäckenområdet
      2 bäckenorgan
      1 bäckenregionen
      1 bäckenreservoar
      1 bäckenringen
      2 bäckenringens
      1 bäckenskål
      1 bäckensnitt
      1 bäckenuppluckring
      1 bäckenutvidgande
      1 backflöde
      1 background
      1 backmark
      1 backronym
      2 backsipporna
      2 backsippssläktet
      1 bäckstränder
      1 backtimjan
      1 backtrav
      1 backventil
      1 bacl
      3 bacon
      1 bacterier
      1 bacteroider
      1 bacteroidetes
      1 bactrim
      1 baculum
     27 bad
     14 bada
    177 båda
      1 badade
      2 bådadera
      1 badande
      1 badanläggningar
      1 badanläggningen
      1 badanläggningens
      5 badar
      1 badaren
      1 badas
      1 badavin
      1 badbehandlingen
      3 bädd
      1 bäddar
      2 baddräkt
      1 baddräkten
      1 baddräktens
      1 bäddvärmare
    473 både
      4 badet
      1 badets
      1 badformer
      4 badger
      2 badhandduk
      9 badhus
      5 badkar
      1 badkarsolyckor
      4 badklåda
      1 badklådan
      1 badkläderna
      1 badkultur
      2 badlakan
      1 badmassagen
      2 badmode
      1 badplatser
      1 badrum
      1 badrummet
      1 badrums
      1 badrumshandduk
      1 badrumsskåp
      1 badstuga
      1 badstugorna
      1 badu
      3 badvakt
      3 badvaktens
      3 badvakter
      1 badvatten
      1 bafucin
      1 bag
      2 bagage
      5 bågar
      2 bagarastma
      1 bagarastmatiker
      1 bägarceller
      1 bägarcellerna
      2 bagare
      2 bägare
      9 bågarna
      1 bägarnattskatta
      1 bågböjda
      1 bågbrillor
      1 bågbrillorna
      1 bagdad
      5 båge
      6 bågen
      1 bågens
      1 bageri
      1 bagg
      1 båggångar
     20 bägge
      2 baggen
      1 baghdad
      1 bågmaterial
      1 bågminuter
      1 bågskytteträning
      1 bågsträngar
      1 bågsträngens
      1 bågsvetsning
      1 baháí
      2 baháíer
      1 baháílitteraturen
      1 baháítron
      1 baháulláhs
      1 bailii
      2 baillie
      2 baillies
      1 bainbridge
      2 bainbridgereflexen
      1 baird
      2 bajonettfattning
      1 bajonettkoppling
      7 bak
      2 bakades
      1 bakar
      2 bakas
     17 bakåt
      1 bakåtböjning
      1 bakåtflödande
      1 bakåtlutande
      1 bakåtneråtrörelser
      1 bakåtriktade
      2 bakben
      2 bakbenen
      1 bakdel
      1 bakelit
      1 bakermanskranenburg
      1 bakfickan
      1 bakfylla
     34 bakgrund
     11 bakgrunden
      1 bakgrundsbullernivån
      1 bakgrundsfärgen
      1 bakgrundsfrekvens
      2 bakgrundsstrålning
      1 bakgrundsstrålningen
      2 bakhåll
      1 bakhållsplats
      1 bakhorn
      2 bakhuvudet
      3 bakifrån
      2 bakkroppen
      2 baklänges
      4 baklob
      1 baklofen
      1 bakluckan
      2 bakning
    102 bakom
     41 bakomliggande
      1 bakomvarande
      1 bakonmliggande
     26 bakre
      4 baksida
      6 baksidan
      1 bakslag
      2 baksmälla
      1 baktassarna
      5 baktericid
      1 baktericida
     41 bakterie
      1 bakterieangrepp
      1 bakterieansamlingar
      1 bakteriearter
      1 bakteriearterna
      1 bakteriebeläggning
      1 bakteriecellens
      2 bakterieceller
      1 bakteriecellerna
      1 bakteriecid
      1 bakteriedna
     14 bakteriedödande
      2 bakteriedysenteri
      6 bakterieflora
      6 bakteriefloran
      1 bakterieförekomst
      1 bakteriefria
      1 bakteriegift
      1 bakteriegifter
      1 bakteriegrupperna
      5 bakterieinfektion
      6 bakterieinfektioner
      1 bakterieinfektionshämmande
      1 bakterieinsjuknandet
      1 bakteriejämvikten
      1 bakteriekänsliga
      1 bakteriekolonier
      1 bakteriekontamination
      2 bakteriekulturer
     69 bakteriell
     15 bakteriella
      1 bakteriellt
      1 bakteriemi
    120 bakterien
     20 bakteriens
      8 bakterieodling
      2 bakterieodlingar
      1 bakterieorsakad
      1 bakterieproteiner
      1 bakterieprov
    321 bakterier
      1 bakterierdet
      1 bakterieresistensen
      1 bakteriergram
      1 bakterierika
     77 bakterierna
      1 bakteriernaclostridium
      7 bakteriernas
      1 bakteriernyttobakerier
      8 bakteriers
      1 bakterieruri
      4 bakteriesjukdom
      1 bakteriesläktet
      3 bakteriestam
      7 bakteriestammar
      1 bakteriestammen
      2 bakteriestammens
      6 bakterietillväxt
      1 bakterietillväxten
      3 bakterietyper
      1 bakterietyperna
      1 bakterieutsatta
      2 bakterieväxt
      1 bakterigruppen
      1 bakteriocidal
      1 bakteriociner
      1 bakteriofagterapi
      3 bakteriologen
      2 bakteriologi
      3 bakteriostatisk
      2 bakteriostatiska
      1 bakteriostatiskt
      1 bakteristammar
      7 bakteriuri
      1 bakterostatiska
      2 baktill
      1 bakvägen
      1 bakväggs
      2 bakvänd
      1 bakvänt
      1 bakverk
      7 bål
      1 balance
      3 balanit
     19 balans
      6 balansen
      1 balansera
      5 balanserad
      3 balanserar
      2 balanseras
      3 balanserat
      2 balansering
      1 balansimpulser
      1 balansnivå
      4 balansorgan
      6 balansorganen
      3 balansorganet
      1 balansövningar
      1 balansrubbningar
      1 balanssinne
      1 balanssinnena
      3 balanssinnet
      1 balansstörningar
      1 balanssvårigheter
      3 balanssystemet
      1 balansteroin
      1 balconette
      2 balconetten
      1 balconnet
      1 baldakiner
      1 balders
     10 bålen
      1 bålens
      1 bålgetingar
      1 balind
      3 balis
      1 balise
      3 balisen
      7 baliser
      5 baliserna
      1 balisfel
      4 balja
      1 baljan
      3 baljkapslar
      2 baljväxter
      1 balkan
      2 balkanhalvön
      1 balkong
      1 ballast
      1 ballistiska
     11 ballong
      1 ballongbrakyterapi
      9 ballongen
      2 ballongkateter
      1 ballongkompression
      1 ballongutvidgningen
      1 ballongvidga
      6 ballongvidgning
      1 bållsjuka
      1 balneoterapi
      1 balsal
      5 balsam
      1 balsambehandling
      1 balsamering
      7 bälte
      4 bältet
      2 baltikum
      1 baltimore
      2 bältor
     23 bältros
      2 bältrosen
      1 bältrosinfektion
      1 balttysk
      1 bälz
      3 bambu
      1 bamburör
      2 ban
      1 bana
      7 banan
      1 banandieten
      2 bananer
      1 bananflugor
      1 banans
      5 banbrytande
      1 banbrytare
      3 bancrofti
     22 band
      3 bandage
      1 bandagebehovet
      1 bandagering
      7 bandbredd
      2 bandbredden
      1 bandbreddsmätning
      3 banden
      4 bandet
      1 bandformiga
      1 banditer
      2 bandler
      3 bandmask
      1 bandmaskarna
      2 bandmått
      2 bandmåttet
      1 bandpassfilter
      1 bands
      1 bandspelarekg
      1 bandunduprovinsen
      1 bandunduregionen
      1 bane
      1 bangalore
      1 bangårdar
      2 bangham
      1 bangladesh
      2 bangs
      2 bank
      3 bänk
      1 bänkar
      1 bänkdiskmaskiner
      3 banken
      1 banker
      1 bankerna
      2 bankkonto
      1 bankkonton
      1 bänkskivor
      1 bannlyst
      1 bannlyste
      1 bano
      3 banor
      1 banorna
      1 bansträcka
      1 bansystemet
      2 banta
      1 bantare
      7 bantaren
      1 bantigenen
      1 bantigenerna
      6 banting
     17 bantning
      2 bantningen
      3 bantningsmedel
      1 bantningsmetoden
      3 bantningsmetoder
      1 bantningspreparat
      1 banvallar
      1 baptiste
     37 bar
      3 bår
     87 bär
    371 bara
     42 bära
      4 bärande
     22 bärare
      8 bäraren
      1 bärarenimmun
      5 bärarens
      1 bärarmolekylen
      1 bärarmolekyler
      2 bärarna
      1 bärarproteinet
      1 bärarskap
     10 bäras
      2 barbae
      3 barbell
      2 barberare
      1 barbershop
      2 barbiturat
      3 barbiturater
      1 barbituraternas
      2 barbro
      3 barbröstade
      1 barcelona
      1 bard
      1 bardot
      1 bardskärare
      1 båren
     17 bären
      1 bärens
      3 barer
      1 bäres
      1 bäret
      3 barfota
      2 barfotaläkare
      1 barfotaläkarna
      1 barfotamedicin
      2 bariatri
      3 bariatrin
      9 barium
      1 bariumförgiftning
      1 bariumhydroxid
      1 bariuminnehållande
      2 bariumjonen
      1 bariumjonerna
      1 bariumklorid
      1 bariumlavemang
      3 bariumnitrat
      2 bariumoxid
      1 bariumsalter
      1 bariumsalterna
      1 bariumsaltförgiftning
     12 bariumsulfat
      1 bariumsulfatets
      2 bariumsulfid
      8 bark
     10 barken
      1 barkley
      1 barkleys
      1 barkliknande
      1 bärliknande
      2 barlind
      1 bärlind
      1 barlinda
      1 barlindemyren
      1 barlow
      1 barmen
    750 barn
      1 barnaåren
      2 barnadödlighet
      4 barnadödligheten
      1 barnadråp
      4 barnafödande
      1 barnaföderskan
      3 barnaföderskor
      1 barnafödsel
      1 barnafödslar
      1 barnamord
      1 barnamordsplakatet
      1 barnanestesin
      1 barnår
      1 barnarbetare
      3 barnarbete
      1 barnard
      3 barnastma
      1 barnavårdscentraler
      1 barnavårdscentralerna
      1 barnbajs
      1 barnbeck
      1 barnbecket
      3 barnbördshus
      1 barnbördshusen
      1 barnbördshuset
      1 barndermatologi
      1 barndet
      1 barndödlighet
      1 barndödligheten
      9 barndom
     29 barndomen
      1 barndomsallergier
      1 barndomsår
      1 barndomsåren
      1 barndomsdöva
      1 barndomstrauma
      1 barndomstrauman
      1 barnemorska
     61 barnen
     10 barnens
      2 barnesi
    194 barnet
     70 barnets
      2 barnfamiljer
      1 barnfänge
      5 barnfetma
      1 barnfetman
      1 barnfobier
      1 barnhälsovård
      1 barnhälsovården
      1 barnhemsbarn
      1 barnhjärtläkare
      1 barnhus
      1 barnkirurgen
      1 barnkirurgi
      7 barnläkare
      6 barnläkaren
      1 barnleksak
      9 barnlöshet
     20 barnmorska
      5 barnmorskan
      2 barnmorskans
      1 barnmorske
      1 barnmorskebok
      1 barnmorskeförbundet
      1 barnmorskegroden
      1 barnmorskemottagning
      1 barnmorskereglemente
      1 barnmorskereglementet
      4 barnmorskeutbildning
      1 barnmorskeutbildningen
      1 barnmorskeyrket
     12 barnmorskor
      7 barnmorskorna
      1 barnmorskornas
      1 barnmottagning
      1 barnmottagningen
      1 barnneurokirurgi
      1 barnomsorgskola
      1 barnortopeder
      1 barnortopedi
      1 barnpsykiater
      1 barnpsykos
      1 barnröst
     17 barns
      3 barnsäng
      1 barnsängen
      2 barnsängens
      6 barnsängsfeber
      4 barnsängsfebern
      2 barnsängsfeberns
      1 barnsängskvinna
      1 barnsängskvinnor
      1 barnsängstiden
      1 barnsbörden
      3 barnsjukdom
      7 barnsjukdomar
      2 barnsjukhus
      1 barnsjukhuset
      1 barnsjukvården
      1 barnsjukvårdens
      1 barnslig
      2 barnspecialist
      1 bärnsten
      1 bärnstenar
      1 barntandborste
      2 barntandkräm
      1 barnuppfostran
      1 barnvaccin
      2 barnvaccination
      1 barnvaccinationerna
      1 barnvaccinationsprogrammet
      1 barnvagn
      1 baron
      1 baroreceptorer
      1 baroreceptorerna
      1 barotramuma
      4 barotrauma
      1 bärplockarsjuka
      3 barr
      1 barrbuske
      6 barren
      1 barrésinoussi
      2 barretts
      6 barriär
      3 barriären
      6 barriärer
      1 barriärfunktion
      1 barriärkräm
      1 barriärmetoder
      1 barriärrevet
      2 barriärskydd
      1 barrier
      1 barrikaderar
      2 barrlind
      2 barrskog
      1 barrskogsplantor
      5 barrträd
      1 barrträds
      2 barrväxt
      1 barrväxterna
      1 barry
      8 bars
     21 bärs
      1 bärsaften
      1 bärsärkagång
      1 bärsärkar
      1 bärsärkaraseri
      1 bärsärkare
      1 barson
      2 bart
      2 bartlett
      1 bartonella
      1 barys
      4 baryt
      1 barytens
     19 bas
      1 basaglia
      2 basal
     14 basala
      1 basalbiologiska
      5 basalcellscancer
      1 basalcellstumör
      1 basaldos
      1 basaldosen
      1 basaliom
      2 basalmembran
      7 basalmembranet
      1 basalomsättning
      2 basalomsättningen
      2 basaltemperatur
      4 basaltemperaturen
      1 basalticus
      1 basartikel
      1 basbehandling
      2 bascentrerat
      2 basel
     10 basen
      4 baser
     15 baserad
     27 baserade
      1 baserades
      6 baserar
     22 baseras
     32 baserat
      1 baserats
      1 basfödan
      1 basform
      1 basfs
      4 basic
      1 basidiesvampar
      3 basilarmembranet
      2 basinsulin
      1 basiron
      4 basis
      2 basisk
      6 basiska
      3 basiskt
      1 baskerna
      2 baskurva
      3 baskurvan
      1 baslinje
      3 baslinjen
      1 basljud
      1 basmedicinska
      1 basmetoden
      1 baso
      1 basofil
      1 basofila
      4 basofiler
      1 basofilerna
      1 basolateralt
      1 baspar
      1 bassängbad
      2 bassängen
      1 bassänger
      1 bassängvatten
      1 bassiasmöret
      2 basspecialitet
      1 basstatens
      2 bast
     69 bäst
     62 bästa
      1 bastarder
      1 bäste
      1 bastet
      1 bastfibrer
      1 bastoner
      1 bastrumman
      1 bästsäljande
      1 bästsäljaren
     17 bastu
      2 bastuaggregatet
      1 bastuaggregatets
      8 bastubad
      2 bastubadandet
      2 bastubadare
      1 bastubadaren
      1 bastubadet
      1 bastubadning
      1 bastuinrättningar
      1 bastuklubbslagen
      1 bastukonstruktionen
      1 bastukultur
      1 bastukvast
      2 bastukvasten
     11 bastun
      1 bastuna
      1 bastuns
      3 bastur
      2 basturuskan
      1 bastutraditionen
      2 bastuträsk
      1 bastuträsket
      1 bastuugn
      1 bastuvärd
      1 basu
      1 basvetenskaplig
      4 båt
      1 bataljonsnivå
      4 båtar
      1 båtars
      1 båthylla
      1 båtlift
      1 båtlika
      2 båtliv
      1 båtlivet
      1 baton
      1 batong
      1 batonger
      1 båts
      3 batson
      8 batteri
      1 batteridriven
      3 batterier
      1 batterierna
      2 batteriet
      1 batteriets
      1 batterimätning
      1 batteritest
      1 batterityp
      2 battista
      1 battle
    179 bättre
      1 bättring
      1 bättringsvägen
      1 bauhin
      1 bauhinii
      1 bauhinska
      1 bausch
      3 bauxit
      1 bäver
      2 bayard
      1 bayer
      1 baylisascariasis
      1 bayliss
      3 bb
      2 bbavdelning
      1 bbavdelningen
      2 bbcs
      2 bbd
      2 bbr
      3 bbrist
      2 bc
      5 bcell
      1 bcellen
     14 bceller
      4 bcellerna
      1 bcellslymfom
      6 bcg
      3 bcgvaccin
      5 bcgvaccinet
      1 bcrabl
      6 bdd
      3 bdelen
      1 bdsm
      1 bdsmsfärerna
     12 be
      1 beach
      1 bead
      1 beaded
      4 beakta
      3 beaktande
      1 beaktar
      1 beaktas
      1 beaktning
      1 bealevägen
      1 bealsio
      8 bearbeta
      4 bearbetad
      1 bearbetades
      5 bearbetar
     11 bearbetas
      1 bearbetat
      2 bearbetats
      7 bearbetning
      2 bearbetningen
      1 bearbetningsareorna
      1 bearbetningsflyt
      1 bearbetningshastighet
      3 beatles
      1 beauterne
      2 bebisens
      1 bebott
      2 bebyggelse
      2 becel
      1 bechterew
      2 bechterews
      1 beck
      1 beckomberga
      1 becl
      1 becquerel
      1 beda
      1 bedlam
     37 bedöma
      1 bedömandet
     11 bedömas
      2 bedömde
      2 bedömdes
     13 bedömer
      1 bedömingslista
     32 bedömning
      8 bedömningar
      1 bedömningarna
     13 bedömningen
      1 bedömningsfråga
      2 bedömningsinstrument
      2 bedömningsnämnden
      1 bedömningsunderlag
      1 bedömningsverktyg
     34 bedöms
      2 bedömt
      4 bedömts
      3 bedöva
      1 bedövad
      1 bedövade
      3 bedövande
      3 bedövar
      3 bedövas
     10 bedövning
     13 bedövningen
      1 bedövningsgasen
      1 bedövningsgel
      7 bedövningsmedel
      1 bedövningsmedlen
      1 bedövningsmedlet
      1 bedövningsplåster
      1 bedövningsspray
      1 bedövningsspruta
      2 bedragare
      1 bedragares
      5 bedrägeri
      1 bedrägerier
      1 bedrägerisituation
      1 bedräglig
      1 bedrägliga
      2 bedrägligt
      2 bedragna
      4 bedrev
      3 bedrevs
      3 bedrift
      2 bedriften
      4 bedriva
      7 bedrivas
     14 bedriver
      3 bedrivit
      4 bedrivits
     38 bedrivs
      1 bedrövande
      1 beduinerna
      1 bee
      1 beersheba
      1 beethoven
      3 befäl
      1 befälen
      1 befälhavare
      2 befälskår
      4 befann
      4 befanns
      1 befarad
      1 befarade
      3 befaras
      1 befarats
      1 befäste
      1 befästningsgördeln
      2 befattning
      1 befattningen
      1 befattningsbenämningen
      2 befattningshavare
      9 befinna
     56 befinner
      5 befintlig
     12 befintliga
      1 befintligt
      2 befogad
      1 befogat
      3 befogenhet
      2 befogenheten
      4 befogenheter
      2 befogenheterna
      2 befolkade
     36 befolkning
      5 befolkningar
      3 befolkningarna
    109 befolkningen
      4 befolkningens
      2 befolknings
      1 befolkningsbegränsning
      1 befolkningsgrupp
      2 befolkningsgrupper
      1 befolkningskontroll
      2 befolkningspolitik
      2 befolkningspolitiken
      1 befolkningspolitikens
      1 befolkningsstatistik
      1 befolkningsstudier
      1 befolkningstalet
      2 befolkningstillväxt
      1 befolkningstryck
      1 befordra
      1 befordran
      1 befordras
      2 before
      1 befrämja
      1 befrämjande
      2 befria
      2 befriad
      1 befriade
      1 befriar
      2 befrias
      1 befriat
      2 befrielse
      8 befrukta
      4 befruktad
     17 befruktade
      1 befruktades
      1 befruktande
      8 befruktar
      7 befruktas
      9 befruktat
     35 befruktning
     20 befruktningen
      1 befruktningsapparat
      2 befruktningsapparaten
      1 befruktningsdugliga
      1 befruktningsorgan
      2 befruktningstillfället
      1 befuktaren
      1 befullmäktigad
      2 befunnit
      5 befunnits
      2 beg
     15 begå
      1 begagna
      1 begagnade
      1 begagnades
      2 begagnat
     17 begår
     13 begär
      7 begära
      2 begäran
      1 begärande
      1 begärde
      2 begäret
      4 begås
     10 begått
      3 begåtts
      1 begav
      1 begåvad
      3 begåvade
     11 begåvning
      1 begåvnings
      1 begåvningsgraden
      1 begåvningshandikapp
      1 begåvningsnivån
      1 begåvningsstödjande
      1 begåvningsstörningar
      1 begåvningsstörningen
      1 begåvningstester
      1 bege
      8 begick
      1 begicks
      1 begränad
     22 begränsa
     50 begränsad
     23 begränsade
      3 begränsades
      4 begränsande
     14 begränsar
     16 begränsas
     23 begränsat
      1 begränsats
      9 begränsning
     18 begränsningar
      1 begränsningarna
      2 begränsningen
      1 begrava
      3 begravas
      1 begravd
      1 begravda
      5 begravning
      1 begravningar
      2 begravningen
      1 begravningsceremonier
      1 begravningsgudstjänst
      1 begravts
     92 begrepp
     18 begreppen
    165 begreppet
      2 begreppets
      2 begreppsbildning
      3 begreppsförvirring
      1 begreppsmässiga
      1 begreppspar
      1 begreppsvärld
      4 begripa
      2 begriplig
      6 begriplighet
      1 begrundan
      1 begs
      4 begynnande
      2 begynnelse
      1 begynnelseljud
      1 begynnelsen
     12 behå
      3 behåar
      3 behåbränning
      1 behäftades
      1 behag
      1 behaga
      1 behagat
      1 behagfulla
      3 behaglig
      1 behagligare
      1 behagligt
      1 behåkupor
      1 behåliknande
      3 behåll
     17 behålla
     17 behållare
      8 behållaren
      1 behållarvärd
      1 behållas
      7 behåller
      3 behållit
      1 behållits
      2 behån
      1 behändigt
    140 behandla
      8 behandlad
     20 behandlade
      8 behandlades
      8 behandlande
     48 behandlar
      3 behandlare
      1 behandlaren
    293 behandlas
      3 behandlat
     15 behandlats
      1 behandligen
    969 behandling
    117 behandlingar
      7 behandlingarna
      1 behandlingarnas
      1 behandlingbart
    298 behandlingen
      4 behandlingens
      1 behandlingform
      1 behandlingkliniker
      1 behandlingmöjligheterna
      1 behandlings
      8 behandlingsalternativ
      2 behandlingsalternativet
      1 behandlingsanläggning
      1 behandlingsåtgärd
      3 behandlingsåtgärder
      1 behandlingsbara
      1 behandlingsbehov
      1 behandlingscykel
      1 behandlingsdilemmat
      2 behandlingseffekt
      2 behandlingsfilosofi
      1 behandlingsförlopp
      2 behandlingsförloppet
     22 behandlingsform
      5 behandlingsformen
     12 behandlingsformer
      1 behandlingsformerna
      1 behandlingsförsök
      5 behandlingshem
      1 behandlingshemmet
      1 behandlingsinsatsen
      2 behandlingsinsatser
      2 behandlingsklinikerna
      2 behandlingskrävande
      1 behandlingskur
      1 behandlingsmål
      1 behandlingsmedel
     18 behandlingsmetod
      7 behandlingsmetoden
     38 behandlingsmetoder
      5 behandlingsmetoderna
      2 behandlingsmöjlighet
      2 behandlingsmöjligheter
      1 behandlingsmöjligheterna
      1 behandlingsområde
      6 behandlingsområdet
      1 behandlingsperioden
      1 behandlingspersonalen
      1 behandlingsplan
      1 behandlingsplanen
      1 behandlingsplanerna
      1 behandlingspremisser
      4 behandlingsprogram
      1 behandlingsregimer
      1 behandlingsregionen
      1 behandlingsrekommendation
      5 behandlingsrekommendationer
      1 behandlingsrekommendationerna
      1 behandlingsrelaterade
      1 behandlingsresistent
      4 behandlingsresultat
      3 behandlingsresultaten
      3 behandlingsresultatet
      1 behandlingsrum
      1 behandlingsrummet
      1 behandlingssätt
      1 behandlingssättet
      3 behandlingsstället
      1 behandlingsstart
      1 behandlingssteget
      1 behandlingsstudier
      1 behandlingssvar
      2 behandlingssvikt
      1 behandlingsteknik
      1 behandlingstekniker
      1 behandlingsterapier
      3 behandlingstid
      4 behandlingstiden
      1 behandlingstider
      1 behandlingstiderna
      1 behandlingstillfälle
      1 behandlingstraditioner
      1 behandlingstypen
      1 behandlingsuppehåll
      1 behandlingsvägar
      2 behandlingsvalet
      1 behandlingsvarianter
      1 behanlingen
      4 behåring
      4 behåringen
      2 behärskar
      1 behavior
      2 behavioral
      1 behaviorism
      1 behaviorismen
      2 behaviorismterapi
      1 behaviorister
      1 behavioristiska
      1 behaviour
      2 behavioural
      2 beh�ets
      2 behjälplig
      1 behjälpligt
      3 behöll
      1 behölls
      1 behörig
      1 behöriga
      8 behörighet
      2 behörigheten
    130 behov
     59 behöva
      3 behövande
     19 behövas
      1 behövd
     16 behövde
      6 behövdes
      4 behoven
    258 behöver
      1 behöves
     23 behovet
      1 behövliga
     98 behövs
      1 behovsbedömning
      2 behovstillfredsställelse
      3 behövt
      2 beige
      1 beigt
      2 being
      1 beir
      4 beivras
      1 bejafolket
      2 bejakas
      3 bejel
      2 bejerot
      1 bejerots
      1 bekämningsmedel
     31 bekämpa
      2 bekämpades
      1 bekämpande
      8 bekämpar
      5 bekämpas
      1 bekämpat
     13 bekämpning
      3 bekämpningen
      1 bekämpningsfrågan
     29 bekämpningsmedel
      4 bekämpningsmedlet
      2 bekämpningsmetoder
      1 bekämpningsprodukter
      1 bekämpningssynpunkt
      1 bekännelse
      3 bekant
      4 bekanta
      1 bekfräftar
      1 beklädd
      1 beklagande
      1 beklämmande
      1 beklätt
      1 bekosta
      1 bekostnad
     14 bekräfta
      2 bekräftad
      7 bekräftade
      3 bekräftades
      3 bekräftande
      3 bekräftar
     13 bekräftas
      2 bekräftat
      6 bekräftats
      4 bekräftelse
      1 bekrigade
      2 bekvämare
      1 bekvämlighetsflagg
      3 bekvämt
      1 bekymmer
      1 bekymrad
      3 belagd
      1 belagda
     20 belägen
      4 beläget
     44 belägg
      1 belägga
      4 beläggas
      2 beläggen
      1 belägger
      6 beläggning
      4 beläggningar
      1 beläggningen
      4 beläggs
      5 belägna
      1 belägrad
      1 belägringen
      5 belagt
      1 belagts
      1 belamring
      1 belamringen
      1 belasta
      1 belästa
      3 belastade
      4 belastar
      1 belastas
     32 belastning
      2 belastningar
     10 belastningen
      1 belastnings
      1 belastningsförmånga
      2 belastningssjukdomarna
      4 belastningsskador
      1 belastningssmärtor
      1 belgian
      7 belgien
      1 belgiens
      4 belgiska
      1 belgiske
      4 bell
      1 bella
      5 belladonna
      1 bellamy
      3 belle
      5 bellman
      3 bells
      1 belönade
      3 belönades
      2 belönande
      1 belönar
      3 belönas
      1 belönats
      5 belöning
      5 belöningar
      2 belöningarna
      1 belöningen
      1 belöningscentra
      1 belöningsrutor
      2 belöningsschema
      1 belöningssystem
      1 belöningssystemet
      1 belopp
      1 below
      1 belphegor
      1 belur
      4 belysa
      2 belysande
      1 belysas
      3 belyser
      2 belyses
      6 belysning
      4 belyst
      1 bemålade
      1 bemannades
      2 bemannas
      1 bemannats
      1 bemanning
      1 bemanningsföretag
     16 bemärkelse
      1 bemärkelsen
      1 bemärkelser
      1 bemästras
      1 bemästringsförmåga
      1 bemödanden
      3 bemöta
      1 bemötabr
      6 bemötande
      1 bemötas
      1 bemöts
      2 bemöttes
    107 ben
      2 bena
      1 benabid
      1 benadanti
      1 benådas
      1 benådats
      3 benägen
     22 benägenhet
      8 benägenheten
      3 benäget
     12 benägna
      2 benämna
      7 benämnas
      5 benämnd
      1 benämnda
      3 benämnde
      6 benämndes
     49 benämning
      9 benämningar
      1 benämningarna
     37 benämningen
     57 benämns
      7 benämnt
      3 benämnts
      2 benandante
     13 benandanti
      1 benandantirättegången
      2 benandantis
      2 benändarna
      1 benbildningen
      1 benbiopsi
      2 benbitar
      1 benbiten
      9 benbrott
      3 benbrytarfeber
      1 bencellerna
      2 bencement
      1 benckiser
      1 bene
      2 benedicks
      1 benedictow
     42 benen
      1 benens
     24 benet
      2 benets
      1 benficka
      1 benfiskar
      2 bengt
      1 benhammare
     15 benhinneinflammation
      1 benhinnorna
      9 benign
     13 benigna
      1 benimplantatet
      1 beninflammation
      1 benjamin
      1 benjamina
      3 benjaminfikus
      2 benjaminfikusen
      1 benkil
      1 benknölen
      1 benknoppar
      1 benmängd
      1 benmängden
      8 benmärg
     23 benmärgen
      2 benmärgens
      1 benmärgscancer
      1 benmärgsceller
      1 benmärgssjukdomar
      2 benmärgssvikt
      5 benmärgstransplantation
      2 benmärgstransplantationer
      1 benmassa
      1 benmaterial
      1 benmatrix
      1 benmineraltätheten
      1 benn
      1 bennedbrytande
      1 bennedbrytning
      1 bennich
      2 bennivå
      1 bennivån
      1 benödem
      1 benpålagringar
      1 benplugg
      2 benproteser
      1 benringen
      1 benröntgen
      2 bensalkoniumklorid
     22 bensår
      1 []bensazepinol
     21 bensen
      3 bensendiol
      1 bensendioler
      1 bensendisulfonsyra
      1 bensenhexafluorid
      1 bensenmolkylen
      1 bensenparadisulfonsyra
      3 bensenring
      3 bensenringar
      1 bensenringen
     14 bensin
      1 bensinbilar
      1 bensindrift
      1 bensinen
      1 bensinfordon
      1 bensinmackar
      1 bensinmotor
      1 bensinmotorer
      1 bensintillsatser
      1 benskivor
      7 benskörhet
      1 benskörheten
      1 benskörhetssjukdomar
      4 bensmärta
      2 bensmärtor
      1 bensoat
     14 bensodiazepiner
      1 bensodiazepinliknande
      1 bensoesyra
      1 bensoesyrans
      2 bensofenon
      3 bensokinon
      3 bensol
      1 bensopyren
      1 bensoylklorid
      4 bensoylperoxid
      1 benstomme
      3 benstommen
      2 benstommens
      1 benstrukturer
      1 benstycke
      1 benstyrka
      2 bensvullnad
      1 bensylalkohol
      1 bensylbensoat
      1 bensylgrupp
      1 bensylpenicillin
      1 bensylsalicylat
      2 bentall
      3 bentäthet
      5 bentätheten
      1 bentäthetsvärde
      1 bentonit
      1 bentoquatam
      1 benvärk
     10 benvävnad
      6 benvävnaden
      1 benvävnadsceller
      1 benvävnadsintegration
      1 benvävnadsligament
      1 benvävsuppmjukning
      1 benvenuto
      1 benzaldehyd
      1 benzatinpenicillin
      2 benzedrine
      1 benzidam
      1 benzimidazolderivat
      1 benzol
      1 beoh
      2 beordrade
      2 beordras
      1 beordrat
      1 bephanten
      3 beprövad
      4 beprövade
      1 beprövas
      1 beprövat
      4 ber
     11 beräkna
      4 beräknad
      4 beräknade
      5 beräknades
      1 beräknande
      9 beräknar
     40 beräknas
      5 beräknat
      5 beräkning
      7 beräkningar
      3 beräkningarna
      4 beräkningen
      1 beräkningsmatriser
      1 beräkningsmetoder
      1 beräkningsprinciperna
      5 berätta
      1 berättade
      1 berättande
     10 berättar
      5 berättas
      1 berättat
      1 berättats
      3 berättelse
      3 berättelsen
      1 berättelsens
      3 berättelser
      1 berättelserna
      5 berättigad
      2 berättigade
      2 berättigar
      1 berberfolket
      4 bereda
      2 beredas
      5 beredd
      1 beredda
      2 bereddes
      1 bereder
     19 beredning
      5 beredningar
      2 beredningen
      5 beredningsform
      2 beredningsformer
      1 beredningsmetod
      1 bereds
      2 beredskap
      1 beredskapsmediciner
      1 bereonde
      2 berett
      1 berfenstam
      4 berg
      1 bergart
      7 bergarter
      1 bergartsbildande
      6 bergen
      1 bergenbelsen
      1 berger
      2 berget
      1 berggrund
      1 berggrunden
      1 bergh
      1 bergig
      1 bergiga
      1 bergkristall
      1 berglind
      1 berglund
      1 berglunds
      1 bergmark
      1 bergmynta
      1 bergsalt
      1 bergsfriden
      2 bergskedjan
      1 bergsklättrare
      1 bergsklättrarna
      1 bergsklättring
      1 bergslagen
      1 bergsområden
      1 bergson
      1 bergsprickor
      1 bergsregioner
      1 bergsskärningar
      1 bergstrakter
      1 bergvallmosläktet
      2 berikande
      1 berikat
      1 berikning
      1 berit
      1 berkeley
      1 berlandieri
      4 berlin
      1 berlinmurens
      1 berlinpapyrusen
      1 bernadotte
      6 bernard
      2 berne
      1 bernes
      1 bernhard
      1 bernhardii
      1 bernoulliprincipen
    155 bero
     24 berodde
    293 beroende
      1 beroendebehandling
      1 beroendeförhållande
      1 beroendeförhållandet
     12 beroendeframkallande
      1 beroendeläkare
      1 beroendemottagningar
      2 beroenden
      2 beroendeproblematik
     10 beroendet
      1 beroendevård
      1 beroendevården
      2 beröm
      5 berömd
      7 berömda
      1 berömde
      2 berömt
    380 beror
     14 berör
      2 beröra
      1 beröras
      8 berörda
      1 berörde
     35 beröring
      1 beröringen
      1 beröringsfri
      1 beröringskänsel
      3 beröringskänslighet
      1 beröringsöm
      3 beröringspunkter
      1 beröringssignalerna
      8 berörs
      2 berört
      1 berörts
      4 berott
      1 berövade
      1 berövats
      1 berry
      1 berrys
      1 bertel
      1 bertheim
      1 bertianus
      1 bertillonklassificeringen
      1 bertrand
      1 berus
      2 berusad
      1 berusande
      1 berusat
      7 berusning
      1 berusningen
      1 berusningssymptom
      1 beryl
      4 beryll
      2 beryllen
      8 beryllium
      1 berylliumframställning
      1 berylliumhydroxid
      1 berylliumhydroxiden
      4 berylliummetall
      1 berylliummineral
      2 berzelius
      1 besådda
      1 besannats
      3 besatt
      2 besatta
      2 besättelseschamanism
      1 besättelsetrans
      2 besatthet
      1 besattheten
      4 besättning
      2 besättningar
      5 besättningen
      1 besättningsmän
      1 besegrad
      1 besegrats
      1 besicles
      1 besigye
      1 besiktning
      2 besitta
      2 besitter
      1 besjälad
      1 besjungits
      2 besk
      1 beska
      2 beskåda
      4 beskaffenhet
      1 beskällaresjuka
      2 beskärning
      1 beskaste
      6 besked
      2 beskedet
      1 beskedlig
      1 beskedligt
      1 beskhet
      1 beskjuta
     37 beskrev
     45 beskrevs
     41 beskriva
      1 beskrivad
      1 beskrivande
     16 beskrivas
      3 beskriven
     64 beskriver
      2 beskrivet
     10 beskrivit
     20 beskrivits
     19 beskrivna
     41 beskrivning
      6 beskrivningar
      2 beskrivningarna
      9 beskrivningen
     57 beskrivs
      3 besksöta
      1 beskt
      2 beskydd
      1 beskyddare
      1 beskyllningar
      1 beskyllts
      1 beslagtagit
      1 beslagtags
     11 besläktad
     15 besläktade
      9 besläktat
      6 beslöt
      1 beslöts
     26 beslut
      8 besluta
     13 beslutade
      1 beslutades
      3 beslutande
      4 beslutar
      3 beslutas
      3 beslutat
      3 besluten
      8 beslutet
      2 beslutsfattande
      1 beslutsfattare
      1 beslutsfattarna
      1 beslutsförmåga
      1 beslutsträd
      1 besmitta
      4 besoar
      1 besoarantilop
      1 besoargetens
      1 besoarhjort
      1 besoarstenar
     14 besök
      6 besöka
      1 besökande
      7 besökare
      1 besökarna
      6 besöker
      4 besöket
      1 besökshund
      1 besökt
      1 besökte
      1 besöktes
      1 bespottar
      1 bespruta
      1 besprutat
      7 besprutning
      1 besseyre
      6 best
     39 bestå
     77 bestående
      3 beställa
      1 beställas
      1 beställd
      1 beställda
      1 beställer
      1 beställningen
      1 beställt
     14 bestämd
     10 bestämda
      3 bestämde
      1 bestämdes
     33 bestämma
      2 bestämmande
      8 bestämmas
      1 bestämmelse
      1 bestämmelsen
      8 bestämmelser
     10 bestämmer
     10 bestämning
     12 bestäms
     10 bestämt
      6 bestånd
      1 bestånden
      1 beståndet
      2 beständighet
      1 beständigpermanent
      3 beständigt
      1 beståndsbildande
      9 beståndsdel
      9 beståndsdelar
      3 beståndsdelarna
      2 beståndsdelen
    329 består
      1 bestått
     11 besten
      2 bestens
      1 bestfoods
      4 bestick
      1 bestigningen
     22 bestod
      1 bestraffa
      2 bestraffade
      1 bestraffande
      3 bestraffas
      4 bestraffning
      2 bestraffningar
      2 bestrålade
      3 bestrålas
      2 bestrålat
      1 bestrålats
      5 bestrålning
      2 bestrålningen
      1 bestrålningens
      1 bestreds
      1 bestrida
      1 bestritt
      1 bestryka
      1 bestulit
      1 besuch
    113 besvär
      2 besvara
      1 besvarad
      1 besvarade
      8 besvärande
      1 besvärar
      2 besvaras
      4 besväras
     38 besvären
      1 besvärjelser
      2 besvärlig
      3 besvärliga
      1 besvärligaste
      6 besvärligt
      1 besvärsfri
      1 besvärsfria
      1 besviken
      2 besynnerliga
      1 besynnerligt
      2 bet
      8 beta
      4 betaagonist
      3 betaagonister
      1 betaamyloid
      1 betablockad
      2 betablockare
      5 betablockerare
      4 betaceller
      1 betäckning
      2 betade
      1 betaflak
      1 betaglukos
      1 betahemolyserande
      2 betahemolytisk
      4 betahemolytiska
     12 betala
      1 betalactamases
      1 betalades
      2 betalaktam
      6 betalaktamantibiotika
      1 betalaktamas
      1 betalaktamasenzymer
      1 betalaktamaser
      1 betalaktamasstabila
      1 betalaktambindningen
      7 betalaktamer
      1 betalaktamresistens
      1 betalaktamringen
      4 betalar
      1 betalare
      1 betalares
      1 betalas
      1 betalat
      1 betald
      3 betalning
      1 betalt
      1 betamax
      2 betande
      2 betänkande
      1 betänkligheter
      1 betaplussönderfall
      1 betapyrinoskonformationen
      4 betar
      1 betareceptorer
      1 betasönderfall
      1 betastimulerare
      1 betastrålning
      7 bete
     13 beteckna
      2 betecknad
      7 betecknade
      1 betecknande
     27 betecknar
     19 betecknas
      1 betecknat
      2 betecknats
     34 beteckning
      1 beteckningar
      1 beteckningarna
     22 beteckningen
      1 beteckningssätt
    113 beteende
      1 betéende
      3 beteendeaktivering
      3 beteendeanalys
      1 beteendeåtgärder
      1 beteendebehandlingen
      1 beteendeekologi
      1 beteendefokuserad
      1 beteendeförändring
      2 beteendeförändringar
      1 beteendeförändringarna
      1 beteendeforskare
      4 beteendeinriktad
      1 beteendemängden
      6 beteendemässiga
      6 beteendemönster
     52 beteenden
      2 beteendena
      1 beteendendena
      2 beteendepsykologiska
      1 beteenderelaterad
      1 beteenderesponser
      1 beteendestörning
      4 beteendestörningar
      1 beteendestörningen
      2 beteendestudier
      1 beteendesvårigheter
      2 beteendesyndrom
     34 beteendet
      1 beteendetekniker
      1 beteendeterapeutisk
      1 beteendeterapeutiska
     38 beteendeterapi
      1 beteendeterapikbt
      2 beteendeterapin
      1 beteendeuttryck
      1 beteendevetenskap
      1 betelnöt
      1 beten
      4 beter
      1 betesdjuren
      1 betesfeber
      1 beteshagar
      1 betinga
     14 betingad
      9 betingade
      1 betingande
      2 betingar
      2 betingas
      3 betingat
      8 betingelser
      3 betingelserna
     16 betingning
      1 betjänats
      1 betjäning
      1 betjänt
      1 betlehem
      1 betning
      3 beto
      8 betona
      4 betonade
      2 betonades
     14 betonar
      4 betonas
      2 betonat
      1 betong
      2 betongen
      1 betoning
      1 betoningar
      1 betoningen
     13 beträffande
      5 beträffar
     21 betrakta
      2 betraktad
      7 betraktade
      9 betraktades
     12 betraktar
      2 betraktaren
      1 betraktarens
     91 betraktas
      2 betraktat
     10 betraktats
      1 bets
     33 bett
      1 bettelheim
      3 betten
      1 better
      6 bettet
      1 bettets
      2 bettfel
      1 bettfysiologi
      4 bettskena
      3 bettskenan
      2 bettskenor
      1 bettstället
      1 betula
      1 betvivla
      1 betvivlas
      2 between
      8 betyda
     38 betydande
      6 betydde
    120 betydelse
      5 betydelsefull
      9 betydelsefulla
      2 betydelsefullt
      1 betydelselös
      1 betydelselösa
     41 betydelsen
      8 betydelser
      1 betydelseskiljande
      1 betydelseutveckling
    186 betyder
      1 betydesefullaste
      2 betydlig
      1 betydliga
    100 betydligt
      4 betyg
      1 betytt
      1 beundrandet
      1 beundrare
      5 bevaka
      2 bevakas
      4 bevakning
     13 bevakningsföretag
      2 bevakningsföretagen
      1 bevakningsföretagenmarknaden
      3 bevakningsföretagens
      1 bevakningsföretaget
      1 bevakningsföretagets
      1 bevakningsmarknaden
      1 bevakningsstyrka
      1 bevakningsteknik
      1 bevakningstjänst
      2 bevakningstjänster
      1 bevakningstjänsterna
      1 bevakningsverksamhet
      1 bevandrad
      1 beväpnad
      1 beväpnat
      6 bevara
      3 bevarad
      6 bevarade
      4 bevarades
      1 bevarandebiologin
      1 bevarandemodell
      3 bevarar
      4 bevaras
      1 bevarat
      1 beväringar
      2 beväxning
      1 bevekelsegrunderna
      1 beverages
      1 bevf
      1 bevilja
      2 beviljad
      1 beviljade
      1 beviljades
      1 beviljar
      5 beviljas
      1 beviljat
      1 beviljats
     45 bevis
      8 bevisa
      4 bevisad
      5 bevisade
      1 bevisades
      1 bevisar
      4 bevisas
      6 bevisat
      7 bevisats
      1 bevisbara
      5 bevisen
      2 beviset
      7 bevisligen
      1 bevisningen
      1 bevittna
      1 bevittnade
      1 bevittnat
      2 bevl
      1 bezalip
      1 bezoar
      1 bezoldjarisch
      1 bf
      1 bfgf
      1 bfs
     15 bh
      1 bhagavadgita
      1 bhairavi
      1 bhajan
      1 bhaktiyoga
      1 bhlösa
      2 bhn
      2 bhns
      1 bhstorlek
      2 bhstorlekar
      1 bhunderklänning
      1 bhv
      3 bi
      1 biafra
      3 bias
      1 biawak
      1 biaxel
     17 bibehålla
      1 bibehållande
      4 bibehållen
      2 bibehåller
      1 bibehållet
      3 bibehållit
      3 bibehålls
      1 bibehöll
      1 bibehölls
      1 bibel
      1 bibelcitat
     10 bibeln
      1 bibelns
      1 bibelverser
      5 bibliotek
      1 bibliotekarie
      2 bibliotekarien
      1 biblioterapeut
      3 biblioterapeutiska
      6 biblioterapi
      7 biblioterapin
      1 biblisk
      1 bicameral
      5 bic�tre
      1 bidé
      1 bidens
      1 bidi
      1 bidning
     45 bidra
     12 bidrag
      1 bidraga
     19 bidragande
      1 bidrager
     15 bidragit
      1 bidragsfusk
      2 bidragsgivare
      1 bidragsgivarna
     54 bidrar
      8 bidrog
      1 bidrottninggelé
      1 bie
      7 bieffekt
      1 bieffekten
     16 bieffekter
      1 bieffekterna
      1 bienner
      1 biennerna
      1 bien�tre
      1 biersack
      3 bifasisk
      2 bifasiska
      2 bifenyler
      3 bifida
      4 bifidobakterier
      4 bifokala
      1 bifölls
      1 bifynd
      2 big
      1 bigetinggift
      2 bihåla
      2 bihålan
     10 bihåleinflammation
      1 bihåleinflammationer
      1 bihåleslemhinnor
      3 bihålespolning
      6 bihålor
      8 bihålorna
      1 bihålornan
      1 bihålornas
      5 bihang
      6 bihanget
      1 bihangets
      1 bijugatus
      1 bikameralt
     11 bikarbonat
      1 bikarbonatjon
      1 bikarbonatjoner
      2 bikini
      1 bikinibandet
      1 bikinibyxa
      1 bikinilinjen
      3 bikinin
      1 bikiniöverdelen
      2 bikinisnitt
      1 bikinitoppar
      1 bikramyoga
      4 bikrona
      1 bikten
      1 bikuspidalklaffen
     14 bil
      2 bilaga
      9 bilar
      2 bilarna
      1 bilars
      4 bilateral
      6 bilaterala
      1 bilateralsymmetriska
      4 bilateralt
      3 bilavgaser
      1 bilbränsle
     54 bild
     92 bilda
      1 bildäck
      1 bildad
      7 bildade
     25 bildades
      3 bildande
     19 bildandet
    174 bildar
    275 bildas
     12 bildat
      1 bildåtergivning
     23 bildats
      1 bildbaserade
      1 bildbehandlar
      1 bildbehandling
      4 bilddiagnostik
      1 bilddiagnostikverktyg
      1 bildelement
     36 bilden
      1 bildens
     35 bilder
     11 bilderna
      1 bildgivande
      2 bildkvalitet
      1 bildkvaliteten
      1 bildlänkarna
      2 bildligt
      1 bildmottagaren
     17 bildning
      6 bildningen
      1 bildningens
      1 bildprogram
      1 bildrören
      1 bildrörets
      1 bildseendet
      7 bildskärm
      2 bildskärmar
      1 bildskärmsarbete
      1 bildskärmssjuka
      2 bildtelefon
      3 bildtelefoner
      2 bildtelefoni
      1 bildtyper
      1 bildupplösning
      1 bildupptagning
      5 bilen
      1 bilfläktar
      1 bilförare
      1 bilhandlaren
      1 bilharz
      3 bilharzia
      2 bilharzios
      1 bilharziosis
      1 biliär
      1 biliaris
      1 bilious
     26 bilirubin
      3 bilirubinet
      1 bilirubinhalter
      1 bilirubinstegring
      1 bilis
      1 biljard
      1 biljoner
      1 biljud
      1 bilkö
      3 bilkörning
      1 bilkrock
      4 bill
      1 billack
      4 billig
      7 billiga
     16 billigare
      1 billigaste
      7 billigt
      1 billingsmetoden
      2 billroth
      2 biloba
      3 bilolycka
      1 bilolyckor
      1 bilresa
      1 bilresor
      1 biltoga
      1 biltrafiken
      1 bim
      7 bin
      2 bina
      1 binära
      2 binärt
      1 binatus
      1 binaurala
     56 binda
      2 bindan
      5 bindande
      4 bindas
      2 bindehinna
      3 bindemedel
     79 binder
      1 bindevävnad
      1 bindhinna
      4 bindhinnan
      1 bindhinneinflammation
      1 bindhinnekatarr
      2 binding
      1 bindingarna
      1 bindingen
      8 bindning
      3 bindningar
      2 �bindningar
      3 bindningen
      1 bindningsställen
      1 bindningsställena
      1 bindningstal
      1 bindningsyta
      9 bindor
      1 bindorna
     12 binds
     27 bindväv
     12 bindväven
      1 bindvävnaden
      1 bindvävsbildning
      1 bindvävsceller
      1 bindvävsfibrer
      1 bindvävsförändring
      1 bindvävshinna
      1 bindvävskapsel
      1 bindvävsökning
      1 bindvävsrum
      1 bindvävssjukdom
      1 bindvävssjukdomar
      1 bindvävstrådar
      1 bindvävstumör
      2 binet
      1 bingen
      1 binges
      1 binjurar
     16 binjurarna
      1 binjurarnas
      2 binjure
      6 binjurebarken
      1 binjurebarkhormoner
      1 binjurebarkshormoner
      1 binjurebarkssvikt
      1 binjurebarkstimulerande
      3 binjuremärgen
      4 binjuren
      1 binokel
      1 binokeln
      2 binokulära
      1 binokulärt
      6 bioackumulation
      1 bioackumulerande
      1 bioackumuleras
      1 bioackumulering
      1 bioaktiva
      1 bioaktivering
      3 biobädd
      1 biobädden
      1 biobränslen
      1 biocid
      3 biocider
      2 biocidprodukter
      2 bioeffects
      1 bioelectromagnetics
      1 bioetanol
      2 biofilm
      1 biofilmmikrobiologisk
      1 bioflavonoider
      1 biofysiskt
      1 biogaia
      1 biogas
      6 biogena
      1 biografer
      1 biograferna
      1 biografi
      1 biografiska
      1 bioimpedansvåg
      1 bioiniativerapporten
      1 bioinitativerapporten
      1 bioinitiative
      1 bioinitiativerapporten
      2 bioinitiatives
      1 bioinitiativrapporten
      6 biokemi
      5 biokemisk
      7 biokemiska
      3 biokemiskt
      2 biokemisten
      1 biokompatibelt
      1 biokompatibilitet
      2 biolog
      1 biologen
      4 biologer
     13 biologi
      3 biological
      1 biologin
      1 biologisera
     36 biologisk
     74 biologiska
      1 biologiskmekanistika
     32 biologiskt
      1 biology
      1 bioluminiscens
      2 biomagnificeras
      2 biomagnifikation
      1 biomarker
      1 biomarkers
      2 biomassa
      1 biomassan
      1 biomassaträ
      5 biomedicinsk
      1 biomedicinska
      4 biomekanik
      1 biomimetiskt
      4 biomolekyler
      1 biopolymerer
     24 biopsi
      3 biopsier
      1 biopsin
      1 biopsitagning
      1 bioresonans
      4 bios
      1 biosalong
      1 biostatiska
      3 biostatistik
      1 biostatistiska
      1 biostimulerande
      3 biosyntes
      2 biosyntesen
      1 bioteknik
      1 bioteknikcenter
      1 bioteknikmetod
      2 bioterrorism
      8 biotillgänglighet
      3 biotillgängligheten
      2 biotin
      1 biotinidasbrist
      1 biotininfärning
      1 biotop
      2 biotoper
      1 biotransformation
      1 biotransformera
      1 biovetenskap
      1 bipacksedel
     18 bipolär
      6 bipolära
      1 bipolärt
     13 biprodukt
      1 bircks
      1 birgisson
      1 birgitta
      1 birka
      1 birkenau
      1 birklandeyes
      1 birot
      1 birth
      1 bisamhället
      1 bisarr
     11 bisarra
      2 bisarrt
      1 bischinger
      1 bisdesmetioxicurcumin
      1 bisexualitet
      1 bisexuell
      2 bisexuella
      1 bisfenol
      1 bisfenoler
      4 bisfosfonater
      1 bisköldkörtlarna
      1 biskop
      2 biskopen
      1 biskopsmössa
      1 biskopsvigning
      1 bison
      1 bisonoxe
      3 bistå
      3 bistånd
      1 bistande
      1 biståndet
      1 biståndsbeslut
      2 biståndshandläggare
      1 biståndshandläggaren
      1 biståndshandläggarna
      4 bistår
      1 bistås
      1 bistod
      1 bistra
     17 bit
      4 bita
      5 bitande
      7 bitar
      1 bitarna
      2 bitas
      3 bitdd
      5 biten
     10 biter
      2 bitestikelinflammation
      2 bitestikeln
      3 bitestiklar
      8 bitestiklarna
      2 bitit
      2 bitits
      1 bitmunstycke
      2 bitna
      1 biträda
      1 biträder
      1 bitransversal
      2 bitrex
      2 bitrörelser
      1 bits
      1 bitsår
      8 bitter
      1 bitterheten
      3 bittermandel
      1 bittermandelolja
      1 bittersalt
      1 bittersöta
      1 bittert
      1 bittervatten
      2 bittra
      1 bituitus
      2 bitvis
      1 bitynien
      1 bivalenta
      2 bivax
     14 biverkan
     22 biverkning
    156 biverkningar
     26 biverkningarna
      2 biverkningen
      1 biverkningsbegreppet
      1 biverkningscentra
      1 biverkningsfri
      3 biverkningsprofil
      1 biverkningsrapport
      1 biverkningsrapporter
      3 biverkningsrapportering
      1 biverkningsreaktion
      1 biverkningsregistret
      1 biverkningsrisken
      1 biverkningsriskerna
      1 biverkningssignaler
      1 bjärt
      1 bjj
      1 bjöds
      6 björk
      2 björkpollen
      1 björkpollenallergiker
      2 björkris
      1 björkruskan
      3 björn
      1 björnfloka
      1 björnskinn
      1 bj�rnebekk
      1 bjursell
      1 bks
     25 bl
     96 bla
     18 blå
      4 blåa
     10 blåaktig
      1 blåbär
      4 black
      2 bläck
      1 bläckfiskar
      1 blackstone
     47 blad
      1 bladätare
      2 bläddra
     48 bladen
      4 bladens
      4 bladet
      4 bladflikar
      2 bladflikarna
      1 bladform
      1 bladformiga
      2 bladgrönsaker
      1 bladguld
      1 bladiga
      1 bladklängen
      2 bladlöss
      1 bladmagen
      1 bladpar
      2 bladparen
      1 bladrosett
      1 bladrosetter
      1 bladsaften
      2 bladskaft
      1 bladskivan
      1 bladslida
      2 bladundersida
      1 bladväxt
      4 bladvecken
      1 blåemaljerad
      3 blåfärgad
      1 blåfärgade
      1 blåfärgat
      2 blåfärgning
      2 blågrå
      1 blågrått
      4 blågrön
      1 blågult
      1 blaiberg
      1 blålila
      7 blåmärke
     14 blåmärken
      1 blåmärket
      1 blåmärksteckning
      1 blånagel
      1 blancfix
   1040 bland
     11 blanda
      4 blandad
      1 bländad
      7 blandade
      2 blandades
      4 blandar
      1 blandare
     38 blandas
      7 blandat
      1 blandats
      1 blandbar
      1 blandbränslen
      1 blandcell
      1 blandförhållandena
      1 blandform
      2 blandformer
      1 blandinkontinens
      1 blandkost
      5 blandmissbruk
      4 blandmissbrukare
     42 blandning
     11 blandningar
      1 blandningarnas
      4 blandningen
      1 blandraser
      1 blandraserna
      1 blandskog
      1 blandskogsvegetation
      1 blankt
      1 blåolja
      1 blåröd
      2 blåröda
     21 blåsa
     19 blåsan
      1 blåsans
      2 blåsas
      1 blåsbeteendet
      2 blåsbildning
      1 blåscancer
      6 blåser
      6 blåses
      4 blåshalskörteln
      1 blåsigt
      2 blåsinstrument
      1 blåsippan
      2 blåsippssläktet
      8 blåskatarr
      2 blåskatarrer
      1 blåskiftande
      1 blåsliknande
      1 blåsljud
      1 blåsmanet
      1 blåsmaneten
      1 blåsmasksjuka
      1 blåsmola
     30 blåsor
      9 blåsorna
      1 blåste
      1 blastkris
      2 blastocyst
      6 blastocysten
      1 blastocyststadiet
      1 blastom
      1 blåstömning
      1 blåstömningsbesvär
      2 blastomyces
      1 blåsträning
      3 blåsvart
      1 blåsvolym
      4 blåsyra
      1 blåsyran
      1 blåtira
      6 blått
      1 blåviolett
      6 blefarit
      1 blefaron
      5 blek
      9 bleka
      2 blekande
      1 blekare
      2 blekas
      1 blekgrönt
      2 blekgula
      2 blekgult
      6 blekhet
      5 blekinge
      1 blekinges
      1 bleklila
     14 blekmedel
      3 blekmedlet
      5 bleknar
      1 bleknat
     15 blekning
      1 blekningar
      1 blekningseffekten
      1 blekningsgel
      1 blekningsmedel
      1 blekningsmedlets
      1 blekpulver
      1 blekröda
      3 bleks
      9 blekt
      1 blektvättvattnet
      1 blekvätska
      1 blekvätskans
      1 blepharicarpus
      9 bleuler
    305 blev
    463 bli
      2 blick
      3 blickar
      5 blicken
      1 blickomfånget
      1 blickpunkt
      1 blickriktning
      1 blickstilla
      1 blidar
      1 blidas
      1 blidka
      1 blifva
      6 blind
     14 blinda
      1 blindas
      1 blindbock
     29 blindhet
      1 blindhetdövhet
      1 blindheten
      2 blindhund
      1 blindskoleläraren
      1 blindskrift
      1 blindspår
      1 blindsportfedrationen
      6 blindtarm
      2 blindtarmar
     13 blindtarmen
      1 blindtarmens
      4 blindtarmsbihanget
      7 blindtarmsinflammation
      1 blindtester
      4 blinka
      5 blinkande
      1 blinkar
      1 blinkning
      2 blinkningar
      2 blinkningsreflexen
      3 blint
    735 blir
      1 bli[r]
      1 bliss
     10 blivande
    208 blivit
      1 blixtljuset
      1 blixtrande
      1 blixtsmärtor
      1 block
      1 blockader
      1 blockämnet
     11 blockera
      1 blockerad
      2 blockerade
     25 blockerar
      9 blockeras
      3 blockerat
      1 blockerats
      5 blockering
      7 blockeringar
      1 blockeringen
      1 blockeringsmedel
    260 blod
     12 blöda
      2 blodådror
      3 blodådrorna
      1 blodämnen
      8 blödande
      7 blödarfeber
      1 blödarsjuk
     11 blödarsjuka
      1 blodätare
      1 blodåterflödet
     13 blodbanan
      2 blodbanor
      3 blodbanorna
      1 blodbehandling
      3 blodbildande
      1 blodbildningen
      1 blodbildningsökande
      3 blodblandad
      1 blodblandat
      1 blodblodkontakt
      1 blodbr
     11 blodbrist
      1 blodburen
      6 blodburna
      5 blodcancer
      1 blodcancerformen
      1 blodcancern
      1 blodcancrar
      1 blodcell
      1 blodcellen
      5 blodceller
      2 blodcellerna
      1 blodcellers
      1 blodcellscancer
      1 blodcellsutveckling
      1 blodcentraler
     11 blodcirkulation
     15 blodcirkulationen
      1 blodcirkulationssystemet
      1 blodcirkulationssytemet
      1 bloddialys
      1 bloddonation
      1 bloddonationer
      1 bloddroppen
      1 blodelektrolyter
      1 bloden
      7 blöder
    397 blodet
     43 blodets
      1 blodfärgad
      6 blodfetter
      1 blodfettsäkande
      1 blodfettshalter
      3 blodfettssänkande
      1 blodfettsvärden
      1 blodfläckar
     13 blodflöde
     37 blodflödet
      1 blodfobi
      2 blodföde
     14 blodförgiftning
      1 blodförgiftningen
      9 blodförlust
      1 blodförlusten
      2 blodförluster
      9 blodförsörjning
      1 blodförsörjningen
      6 blodförtunnande
      1 blodfyllas
      2 blodfylls
      1 blodgasernas
      1 blodgasprov
      1 blodgenomströmning
      2 blodgenomströmningen
      1 blodgivarbuss
      1 blodgivarbussen
      9 blodgivare
      2 blodgivaren
      1 blodgivarkompensation
      2 blodgivarna
      7 blodgivning
      3 blodglukos
      1 blodglukoshalten
      1 blodglukosmätningar
     10 blodgrupp
      2 blodgrupper
      1 blodgruppering
      2 blodgrupperna
      1 blodgruppernas
      2 blodgruppsantigener
      3 blodgruppsdieten
      6 blodgruppssystem
      1 blodgruppstillhörighet
      4 blodhjärnbarriär
     31 blodhjärnbarriären
      1 blod�hjärnbarriären
      5 blodhjärnbarriärens
      1 blodhundar
      1 blodi
     13 blodig
     12 blodiga
      3 blodigel
      6 blodigeln
      1 blodigelns
      1 blödighet
      5 blodiglar
      1 blodigt
      1 blodinfektion
      3 blodinjektionskada
      1 blodkaliumlösning
      1 blodkällan
     97 blodkärl
     37 blodkärlen
      3 blodkärlens
      2 blodkärlet
      1 blodkärlsflätan
      1 blodkärlsinflammation
      1 blodkärlsnybildning
      1 blodkärlsnybildningen
      2 blodkärlsväggarna
      2 blodkärlsväggen
      1 blodkärlsväggens
      1 blodkoagel
      4 blodkoagulation
      5 blodkoagulering
      8 blodkoaguleringen
      1 blodkomponenter
      1 blodkorv
      1 blodkräkning
      5 blodkropp
     89 blodkroppar
      1 blodkropparkommer
     31 blodkropparna
      5 blodkropparnas
      2 blodkroppars
      1 blodkroppen
      1 blodkroppsbildande
      1 blodkroppsmängden
      2 blodkroppsräkning
      1 blodkroppssönderfallet
      1 blodleverans
      1 blodlevrar
      1 blodlevringen
      2 blodmängden
      1 blodmat
      1 blodmatad
      1 blodnedbrytning
     58 blödning
     69 blödningar
      1 blödningarna
      1 blödningarnas
     14 blödningen
      5 blödningens
      2 blödningsbenägenhet
      1 blödningsbenägenheten
      3 blödningsrisk
      3 blödningsrisken
      2 blödningsrubbningar
      1 blödningsstörningar
      1 blödningstendens
      1 blödningstid
      2 blodnivåer
      1 blodnivåerna
      1 blododling
      1 blododlingar
      6 blodomlopp
     37 blodomloppet
      1 blodomloppets
      2 blodöra
      1 blodört
      1 blodörtssläktet
      7 blodpest
     10 blodplasma
      4 blodplasman
      1 blodplasmavolym
     18 blodplättar
      4 blodplättarna
      2 blodplättarnas
      4 blodprodukter
     42 blodpropp
     22 blodproppar
      5 blodproppen
      1 blodproppshämmande
      1 blodproppslösande
      1 blodproteiner
      2 blodproteinet
     30 blodprov
      1 blodproven
     20 blodprover
      4 blodprovet
      3 blodprovstagning
      1 blodprovstagningar
      2 blodprovstester
      1 blodprovsvärden
      1 blodpudding
      1 blodrenande
      1 blodrester
      1 blodröd
      1 blods
      2 blodsband
      1 blodscener
      2 blodserum
      7 blodsjukdomar
      1 blodskam
      3 blödskinn
      3 blodsmitta
     10 blodsocker
      2 blodsockerfall
      3 blodsockerhalt
      5 blodsockerhalten
      1 blodsockerhöjande
      1 blodsockerkontroll
      6 blodsockermätare
      1 blodsockermätning
      3 blodsockernivå
      2 blodsockernivåer
      3 blodsockernivåerna
      8 blodsockernivån
      2 blodsockerreglerande
      1 blodsockerreglering
      1 blodsockersänkande
      1 blodsockervärde
      9 blodsockret
      2 blodsockrets
      2 blodsputum
      1 blodstämmare
      1 blodstämning
      2 blodstatus
      1 blodstimulerande
      1 blodstockning
      1 blodstoppande
      2 blodstörtning
      3 blodströmmen
      6 blodsugande
      1 blodsugare
      1 blodsystemet
      3 blodtest
      5 blodtester
      1 blodtesterna
      1 blodtillflöde
      4 blodtillförsel
      3 blodtillförseln
      6 blodtransfusion
      1 blodtransfusionen
      1 blodtransfusionens
     17 blodtransfusioner
     93 blodtryck
     35 blodtrycket
      1 blodtrycks
      1 blodtrycksbehandling
      7 blodtrycksfall
      1 blodtrycksfallet
      1 blodtryckshöjande
      1 blodtryckskontroller
      1 blodtrycksläkemedel
      3 blodtrycksmanschett
      3 blodtrycksmätning
      2 blodtrycksmediciner
      1 blodtrycksmodifierande
      3 blodtryckssänkande
      2 blodtryckssänkning
      1 blodtrycksstegring
      1 blodutbyte
      1 blodvaggor
      1 blodvaggorna
      1 blodvallningar
      1 blodvärdar
      2 blodvärde
      4 blodvärden
      2 blodvärdena
      2 blodverksamhet
      8 blodvolym
      5 blodvolymen
      3 bloggar
      4 blöja
      1 blöjeksem
      1 blöjor
      1 blom
      1 blombladskransarna
      1 blomfärg
      1 blomflockar
      1 blomkål
      1 blomkålsöron
      1 blomklasar
      2 blomklasarna
      1 blomklasen
      1 blomknopparna
      1 blomkrona
      1 blomkronan
      1 blomkruka
     14 blomma
     14 blomman
      5 blommande
      4 blommans
     31 blommar
      2 blommat
     58 blommor
     38 blommorna
      1 blommornas
      5 blomning
      7 blomningen
      2 blomningstid
      2 blomningstiden
      1 blompip
      1 blompipen
      1 blomsaften
      1 blomsamlingar
      2 blomställningar
      6 blomställningarna
      1 blomstängeln
      1 blomsterbotten
      1 blomsterhandeln
      1 blomsterhuvudena
      1 blomsterkrans
      3 blomsterur
      1 blomstrande
      1 blomstren
      1 blomvatten
      1 blomväxter
      1 blomväxterna
      1 blomväxters
      1 blonda
      1 blonder
      1 blont
      3 blood
      1 blooms
      1 blossa
      1 blossade
      1 blossande
      1 blossar
      1 blosset
      4 blöt
      6 blöta
      1 blötas
      2 blötdjur
      1 blötlagda
      1 blötläggas
      1 blötlägger
      1 blötläggning
      1 blötläggs
      1 blöts
      1 blott
      1 blött
      5 blotta
      1 blötta
      2 blottade
      1 blottande
      1 blottar
      1 blottas
      1 blottats
      1 blotters
      1 blottlagda
      3 blt
      2 blue
      1 blues
      1 bluff
      1 bluffmakare
      1 blundandes
      1 blundar
      1 blundell
     35 bly
      1 blyacetatlösning
      1 blyånga
      1 blyanvändningen
      1 blybaserade
      1 blyförgiftad
      8 blyförgiftning
      1 blyframställning
      1 blyfyllningar
      2 blyg
      2 blygd
      1 blygdben
      1 blygdbenen
      4 blygdbenet
      1 blygdbensfog
      1 blygden
      3 blygdfogen
     10 blygdläpparna
      1 blygdläpparnas
      2 blyghet
      1 blyglete
      2 blygsam
      2 blygsel
      2 blyhaltig
      2 blymalm
      1 blymalmen
      2 blymetall
      9 blymfocyter
      1 blymfocyterna
      2 blymönja
      1 blyoxid
      1 blyplattor
      1 blyreduktionen
      1 blysalter
      1 blysocker
      1 blyte
      1 blytillsats
      2 blyvitt
      1 bma
      2 bmeningokocker
     22 bmi
      1 bmikilogrammeter
      1 bminnesceller
      3 bmj
      1 bmode
      3 bnp
     11 bo
      1 board
      1 boarda
      3 bob
      1 boc
      7 bocavirus
      1 bocavirusen
      1 bocavirusens
      1 bocaviruset
      1 bocavirusethbov
     35 böcker
      4 böckerna
      1 böckers
      3 bod
      2 bodamer
      2 bodbelastning
      2 bodbelastningen
      2 bodde
      1 boden
      1 bodies
      4 bodm�
      4 body
      1 bodyform
      1 bodywork
      1 boehringer
     16 boende
      1 boendeformerna
      1 boerhaave
      2 boet
      1 bofast
      1 bogart
      1 bögcancer
      1 bogors
      1 boh
      1 bohemen
      2 bohr
      3 bohreffekten
      1 bohus
      1 bohuskusten
      6 bohuslän
      1 boikapslar
      1 boissieri
      1 böj
      8 böja
      1 böjbara
      1 böjbart
     10 böjd
      5 böjda
      2 böjen
      3 böjer
      1 böjerruller
      2 böjlig
      3 böjligt
      1 böjning
      2 böjningar
      5 böjs
      1 böjsenor
      1 böjt
      1 böjtplanrekonstruktion
      1 böjveckseksem
     34 bok
      1 boka
      1 bökade
      1 bokas
     20 boken
      1 bokförläggare
      1 bokform
      1 bokhandelsbiträdet
      1 boklusen
      1 bokmärken
      1 boksidor
      1 bokslutet
      9 bokstav
      7 bokstaven
      4 bokstäver
     12 bokstäverna
      1 bokstavlig
      3 bokstavligen
      2 bokstavligt
      1 bokstavsbeteckningar
      1 bokstavsdiagnos
      1 bokstavsvis
      1 bokstavsvisa
      1 boktryckarkonsten
      1 bolag
      1 böld
      8 bölder
      4 bölderna
     13 böldpest
      1 böldskärning
      1 boletaceae
      1 boletus
      2 boliden
      3 böljande
      3 boll
      1 bollar
      1 bollarna
      1 bollkastning
      1 bollträffar
      1 bolm
      1 bolma
      4 bolmört
      2 bolmörten
      1 bolmörtsskivling
      3 bolmörtsskivlingen
      2 bologna
      1 bolognamodellen
      1 bolognastenar
      1 bolognasystemet
      1 bolus
      1 bolusdos
      2 bolzano
      1 bom
      1 bomb
      1 bombades
      1 bombarderbaggen
      1 bombastus
      1 bombay
      2 bomber
      1 bombs
      1 bombshell
      1 bombshellbh
      1 bombshellbhar
      1 bombykol
      5 bommar
      1 bommarna
     17 bomull
      1 bomulls
      1 bomullsbönder
      1 bomullsfrö
      1 bomullsfrotté
      1 bomullshalsduken
      1 bomullshandduk
      1 bomullsodlingar
      2 bomullspinnar
      1 bomullsproduktion
      1 bomullsskörd
      1 bomullstråd
      3 bomullstussar
      5 bon
      5 bön
      1 bona
      1 bonader
      1 bond
      1 bondebefolkningen
      1 bonden
      5 bönder
      2 bönderna
      1 böndernas
      1 bondeståndet
      1 bondeuppror
      1 bondfilmer
      2 bondgård
      1 bondgårdar
      1 bondgårdens
      1 bondsk
      1 bonebreak
      1 böner
      1 bönestunder
      1 bonfanti
      1 bönformad
      1 bong
      2 boning
      1 bönlika
      1 bonnet
      1 bonoplex
      9 bönor
      1 bönorbönprodukter
      1 book
      1 books
      6 boom
      2 boomers
      3 boostbehandling
      1 boottopfärg
      1 boplatser
     18 bor
    353 bör
      1 borago
      1 borax
      1 boraxsyra
      1 borborygmus
      4 bord
      1 börd
      4 börda
      3 bördan
     26 borde
      1 bordeller
      7 borderline
      1 borderlinepersonlighetsstörning
      1 borderlinepsykos
      1 bordet
      6 bordetella
      1 bordetellaarterna
      1 bördiga
      1 bordsautoklaver
      4 bordssalt
      1 bordsytor
      1 borgar
      2 borgarna
      1 borgerskapet
      1 borgerskapets
     57 börja
    149 började
      1 börjades
    199 början
    198 börjar
     45 börjat
      1 born
      1 borna
      3 bornasjuka
      1 bornaviridae
      2 bornavirus
      1 bornaviruset
      1 borneo
      1 bornm
      1 borno
      1 boroxid
      1 borr
      5 borra
      1 borrade
      4 borrar
      1 borrarna
      1 borrat
     33 borrelia
      1 borreliaartrit
      1 borreliabakterien
      2 borreliabakterier
      2 borreliafall
      3 borreliainfektion
      1 borreliainfektionen
      1 borreliainfektioner
      1 borreliarelaterade
      1 borreliaring
      1 borreliasmitta
      1 borreliatesternas
      4 borrelios
      1 borret
      1 borrhål
      1 borrmaskin
      1 borro
      1 borrproceduren
      1 borrvreden
      5 borst
      4 borsta
      4 borstar
      1 borstas
      5 borste
      1 borstens
      2 borsthuvud
      1 borsthuvuden
      1 borstmögel
      4 borstning
      1 borstningstid
      1 borstresultat
      1 borstskador
      1 borststrån
      1 borststråna
      1 borsttvätt
      1 börsvärlden
      6 borsyra
    275 bort
     24 borta
      1 bortanför
      3 bortåt
      1 bortborrade
      1 bortbytingar
      9 bortfall
      1 bortfallen
      2 bortfaller
      1 bortfallet
      2 bortfallssymptom
      1 bortförande
      1 bortförklara
      1 bortförs
      1 bortförsel
      3 bortgång
      1 bortknytning
      1 bortkopplad
      1 bortmätning
      6 bortom
      2 bortoperation
      1 bortopererad
      1 bortopererade
      1 bortopereras
      3 bortopererat
      1 bortopererats
      2 borträknat
      1 bortrensning
      1 bortsatta
      2 bortsättning
      3 bortse
      7 bortsett
      1 bortstötandet
      2 bortstötning
     12 borttagande
      2 borttagandet
      1 borttager
      1 borttaget
      3 borttagna
      7 borttagning
      1 borttogs
      1 bortträngning
      3 bosatt
      1 bosätter
      1 boscalid
      2 bosch
      6 boskap
      1 boskapen
      1 boskapens
      1 boskaps
      1 boskapsbesättningar
      3 boskapspest
      1 boskapspestvirus
      1 boskapssektorn
      1 boskapsskötsel
      6 bosman
      1 bosmandomen
      1 bosört
      1 bosson
      4 bostad
      7 bostaden
      8 bostäder
      1 bostadsanpassning
      1 bostadsanpassningsbidrag
      1 bostadshus
      1 bostadshusen
      1 bostadskö
      1 bostadslösa
      1 bostadsmiljö
      1 bostadsområden
      1 bostadsort
      1 bostadsrätter
      1 bostadsrum
      4 boston
      1 bostonkorsettens
      1 bostonskolan
      9 bot
     59 bota
      1 böta
      9 botad
     10 botade
      1 botades
     13 botande
      1 botanik
      1 botaniker
      2 botanikern
      1 botanisk
      4 botaniska
      1 botaniskt
      1 botany
     12 botar
     21 botas
      1 botat
      3 botats
      1 botbar
      1 botbara
      1 botbart
     23 botemedel
      1 botemedlet
      1 botemetod
      1 botemetoder
      2 boten
     12 böter
      1 bötfälldes
      2 botgörartåg
      3 botgöring
      1 bothrops
      1 botningsbara
      2 botox
      2 botoxinjektioner
      3 botrytis
      1 bott
      8 botten
      6 bottenfärg
      2 bottenfärgen
      1 bottenfärger
      1 bottensediment
      1 bottenslammet
      2 bottenvåningen
      5 bottnar
      3 bottnen
      7 botulinum
      2 botulinumbakterien
      1 botulinumförgiftning
     10 botulinumtoxin
      1 botulinumtoxinet
      1 botulinustoxin
      4 botulism
      1 botulus
      1 bouchardat
      2 boudin
      2 bourgeois
      2 boven
      2 boverket
      3 bovete
      1 bovin
      2 bovine
      4 bovis
      3 bowl
     11 bowlby
      4 bowlbys
      1 bowles
      1 boxaren
      4 boxning
      1 boy
      1 boyes
      2 boyles
      1 boys
      1 bp
      1 bpatienter
      1 bpositiva
      2 bprs
      5 bqm
      2 bqm�
      1 bqtimmarm
     51 br
    174 bra
      1 brachialis
      1 brachycalyx
      1 brachycephal
      1 brachypterus
      2 brachys
      4 brachyterapi
     15 bråck
      2 bråckbildning
      8 bråcket
      2 brackets
      2 bråckets
      1 bräckliga
      1 bråckliknande
      1 bråcksäck
      1 bråcksäcken
      1 bråckstället
      1 bracteata
      1 brad
      1 bräda
      1 bradbury
      1 brådska
      2 brådskande
      4 bradykardi
      3 bradykinin
      1 bradytakysyndrom
      1 bradytakysyndromet
      1 bradyzoiter
      1 bragte
      4 brahman
      1 braille
      1 braillebokstäverna
      1 brailleskrift
      6 brain
      1 brainbow
      1 brainstorming
      1 braithwaite
      1 bråk
      1 bräkande
      1 brakare
      2 bråkdel
      1 brakfis
      1 bråkiga
      1 brakskit
      1 brakycefal
     71 brakyterapi
      1 brakyterapiingrepp
      1 brakyterapikälla
      2 brakyterapimetoder
      2 brakyterapin
      2 brakyterapins
      1 bräm
      1 branca
      1 branchingenzym
      8 brand
      3 bränd
      1 brända
      1 brandbekämpning
      1 brandbilar
      3 brände
      1 branden
      5 bränder
      1 bränderna
      3 brändes
      1 brandfarlig
      1 brandfarligt
      1 brandgul
      2 brandmän
      1 brando
      1 brandrelaterade
      1 brandröksförgiftning
      2 brandskydd
      1 brandskyddande
      1 brandskyddsmaterial
      1 brandsläckande
      1 brandsläckning
      1 brandsläckningsmaterial
      3 brandt
      1 brandtåligt
      2 brandy
      2 brånemark
      2 brånemarks
      8 bränna
     14 brännande
      1 brännas
      3 brännässla
      2 brännässlan
      1 brännässlans
      2 brännässlor
      2 brännbara
      2 brännbart
      6 bränner
      2 brännhår
      1 bränning
      1 brännmanet
      1 brännmaneterna
      9 bränns
      8 brännsår
      9 brännskada
      2 brännskadad
      1 brännskadade
      5 brännskadan
      1 brännskadas
      1 brännskadats
      1 brännskadeliknande
      1 brännskadevård
     27 brännskador
      1 brännvidder
      1 brännvidderna
      1 brännvin
      1 brännvinskrydda
      2 bransch
      2 branschen
      1 branscher
      1 branschorganisation
      2 branschorganisationen
      8 bränsle
      1 bränsleenergi
      2 bränsleförbrukningen
      1 bränslen
      1 bränslet
      1 bränslevärde
      2 brant
      1 bränt
      1 branta
      1 brantare
      1 branting
      1 brantly
      2 bränts
      2 brasiliansk
      3 brasilianska
     18 brasilien
      1 bråska
      2 brässen
      1 brassicae
      1 brassi�re
      1 brassi�res
      3 bratman
      1 bråttom
      1 braun
      1 brblodet
      3 brbr
      2 brca
      3 breakbone
      1 breakdown
      1 breakheart
      1 breasts
     22 bred
     21 breda
      9 bredare
      1 bredast
      1 bredbands
      1 bredbandsuppkoppling
      6 bredd
      2 bredda
      1 breddas
      4 bredden
      1 breddökat
      2 breder
      1 bredsida
      1 bredspektrigt
      4 bredspektrumantibiotika
      1 bredspektrumantibiotikum
      2 bredspektrumpenicilliner
     10 bredvid
      4 brehmer
      1 bremsstrahlung
      1 brené
      1 brenligt
      1 bresiljaextrakt
      1 breslau
     24 brett
      1 brettanomyces
      6 brev
      1 breven
      1 brevet
      1 brevifolia
      1 brevlådan
      1 brevoxyl
      1 brevromanen
      1 breyers
      1 brföräldraföreningen
      1 brhattrayi
      1 br�hmaa
      2 brian
      1 bricanyl
      1 brider
      1 brides
      2 bridreaktorer
      1 bridreaktorteknologi
      2 brief
      1 brieger
      1 bright
      1 brights
      1 brigitte
      1 brilla
      1 brillenhematom
      2 brillor
      1 brillorna
      2 bringa
      1 bringas
      1 bringats
      3 brinna
      6 brinnande
      8 brinner
      1 brip
    120 brist
      2 brista
     39 bristande
      1 bristel
      1 bristelborste
      2 bristelborsten
     13 bristen
     40 brister
      2 bristerna
     11 bristfällig
      2 bristfälliga
      1 bristfälligt
     11 bristningar
      1 bristningarna
      1 bristningen
      2 bristolmyers
      3 bristsjukdom
      4 bristsjukdomar
      1 bristsjukdomarna
      1 bristsjukdomen
      2 bristsymptom
      3 bristtillstånd
      1 britannien
      9 british
      2 brits
      1 britt
      1 britten
      1 britterna
      7 brittisk
     20 brittiska
      5 brittiske
      1 brittisknederländskt
      2 brittiskt
      1 briva
      3 bro
      1 broad
      3 broar
      4 brocas
      3 broccoli
      7 bröd
      2 broder
      1 broderat
      2 broderier
      1 brodern
      1 broderskap
      2 brodmannarea
      1 brodmannareorna
      1 brödransoner
      1 brody
      1 brokbladig
      1 brokiga
      2 bröllop
      3 brom
      1 bromanders
      1 bromatom
      1 brometan
      1 bromfenoler
      1 bromid
      2 bromiden
      1 bromider
      1 bromintag
      2 bromism
      1 bromismen
      4 brommetan
      5 bromoform
      8 bromsa
      1 bromsade
      5 bromsar
      1 bromsarna
      4 bromsas
      1 bromsbackar
      1 bromsband
      1 bromsbandsfabriken
      1 bromsbelägg
      2 bromsdetaljer
      1 bromshandtag
      1 bromsklossar
      5 bromsljus
      5 bromsmediciner
      1 bromsmedicinerna
      1 bromsmediciners
      2 bromssträckan
      2 bromsstrålning
      1 bromsstrålningen
      1 bromsvätska
      1 bromvatten
      1 bron
      1 bronchiale
      1 bronchiolitis
      4 bronchiseptica
      1 bronchispetica
      3 bronfort
      1 bronk
      1 bronkektasier
      1 bronkepitelet
      2 bronker
      5 bronkerna
      2 bronkernas
      1 bronki
      1 bronkialandning
      1 bronkialastma
      1 bronkialcancer
      1 bronkialmusklerna
      1 bronkialprovokation
      2 bronkiektasi
      2 bronkiektasier
      1 bronkiell
      1 bronkiella
      3 bronkioler
      4 bronkiolerna
      9 bronkiolit
      1 bronkiolitassocierad
      5 bronkit
      7 bronkkonstriktion
      2 bronkopneumoni
      1 bronkopulmunär
      2 bronkoskop
      3 bronkoskopet
      3 bronkoskopi
      1 bronkoskopin
      1 bronkoskopiundersökning
      2 bronkospasm
      1 bronkospasmsymtom
      1 bronkväggen
      4 brons
      2 bronsålder
      4 bronsåldern
      1 bronsåldersrudiment
      2 bronstein
      1 brooke
      2 brooklyn
      1 brookscole
      1 broöppningen
      1 bropelare
      2 bror
      2 broschyrerna
     12 brosk
      1 broskartat
      1 broskdelar
      1 broskdelen
      1 brosken
      5 brosket
      1 broskfisk
      1 broskfiskar
      1 broskflik
      1 broskfogar
      2 broskfogarna
      1 brosksegment
      1 broskstruktur
      2 broskvävnad
     63 bröst
      1 bröståkomma
      1 bröstavledning
      2 bröstavledningar
      2 bröstavledningarna
      2 bröstben
      9 bröstbenet
      1 bröstbestrålning
      1 bröstbesvär
      2 bröstbevarande
      1 bröstbinda
     89 bröstcancer
      1 bröstcancermedicinerna
      1 bröstcancermetastas
      1 bröstcancerpatienter
      1 bröstcancervarianter
      1 bröstcancrar
     58 brösten
      5 bröstens
     58 bröstet
      2 bröstets
      1 bröstfetischism
      1 bröstfickan
      6 bröstfixering
      1 bröstförminskande
      4 bröstförminskning
      1 bröstförminskningskirurgi
      3 bröstförstoring
      1 brösthålan
      1 brösthållare
      2 brösthållaren
      1 brösthälsovården
      1 brösthypertrofi
      8 bröstimplantat
      1 bröstinflammation
      1 bröstkirurgi
      1 bröstkompression
      7 bröstkorg
     31 bröstkorgen
      5 bröstkorgens
      2 bröstkorgsväggen
      1 bröstkörtel
      1 bröstkörteln
      1 bröstkörtelvävnaden
      4 bröstkörtlar
     10 bröstkörtlarna
      1 bröstlapp
      1 bröstlappar
      2 bröstmassa
      2 bröstmassan
     15 bröstmjölk
      1 bröstmjölken
      2 bröstmjölksutsöndring
      1 bröstmjölkutsöndringen
      2 bröstmuskeln
      1 bröstmusklerna
      1 bröstolja
      1 bröstoperationer
      3 bröstpump
      1 bröstpumpen
      2 bröstreduktion
      1 bröstreduktioner
      1 bröstrustningar
      1 bröstrustningarna
      1 bröstsegment
      1 bröstsjukdomar
      7 bröstsmärta
      6 bröstsmärtor
      1 bröstsnörning
      1 bröststorlek
      5 bröststorleken
      2 bröstsymtom
      1 brösttillväxt
      1 brösttumörer
      2 bröstutveckling
      5 bröstutvecklingen
      2 bröstväggen
      4 bröstvårta
     16 bröstvårtan
      6 bröstvårtor
     13 bröstvårtorna
      1 bröstvårtspiercing
     10 bröstvävnad
      4 bröstvävnaden
      1 brösvävnad
      9 bröt
      4 brothers
      3 bröts
     62 brott
      1 brottaröron
      2 brottas
      1 brottens
      9 brottet
      1 brottets
      1 brottmål
      1 brottmålsdomstolen
      3 brottning
      1 brottningsmattan
      1 brottsbalken
      1 brottsbekämpande
      2 brottsbekämpning
      1 brottsförebyggande
      2 brottslig
      3 brottsliga
      8 brottslighet
      2 brottsligheten
      1 brottslighetens
      1 brottsligt
      3 brottsling
      2 brottslingar
      4 brottslingen
      1 brottsoffer
      1 brottsoffren
      2 brottsplatsundersökningar
      1 brottsrubricering
      1 brottstället
      1 brottsteknik
      1 brottsteknikerna
      1 brottstyp
      2 brottsutredning
      1 brottytan
      1 brown
      1 browning
      1 brstorbritannien
      1 brsvenska
      1 bruce
      5 brucei
      1 brucellos
      1 bruch
      2 brucin
      2 brudkrona
      1 brudkronor
      1 brudnäsduken
      3 brudzinskis
      3 brugia
     70 bruk
      4 bruka
     14 brukade
      5 brukades
    323 brukar
      1 brukardrivna
      6 brukare
      3 brukaren
      2 brukarländerna
      1 brukarleden
      1 brukars
      7 brukas
      2 brukat
      3 brukats
     13 bruket
      1 brukettekniken
      1 brukligt
      1 bruksgården
      1 bruksorten
      1 bruksvara
     13 brun
      7 bruna
      3 brunaktig
      2 brunbjörn
      1 brunfärgad
      1 brunfärgat
      1 brungul
      2 brunlila
      5 brunnar
      1 brunnit
      1 bruno
      1 brunögd
      1 brunolivgrön
      1 brunråttan
      1 brunrosa
      1 brunrött
      1 brunstcykel
      1 brunster
      2 brunstighet
      1 brunsvart
      7 brunt
      6 brus
      1 brusande
      1 brusreduktion
      1 brussignaler
      1 brustabletter
      1 brusten
      2 brustet
      1 brustit
      2 brustna
      1 brutala
      2 bruten
      7 brutit
      7 brutits
      2 brutna
      1 bruxellensis
      4 bruxism
      1 bruxismen
      2 bry
      3 bryan
      1 brydestuga
      1 brygd
      1 brygga
      1 bryggor
      1 bryggs
      1 bryn
      1 bryning
      1 bryningen
      3 bryonia
      1 bryophyllum
      4 bryr
     45 bryta
     15 brytas
     65 bryter
      3 brytkraft
      1 brytkraften
      4 brytning
      3 brytningsfel
      2 brytningsfelet
      2 brytningsindex
     57 bryts
      1 brytvärda
      3 bsc
      3 bse
      1 bsefria
      1 bsl
      5 bstreptokocker
      1 bstreptokockinfektioner
      1 bsymtom
      1 bta
      1 b�te
      1 bti
      1 btyp
      1 bu
      1 buaja
      1 bubbelbad
      1 bubbelbildning
      1 bubbla
      1 bubblande
      2 bubblas
      8 bubblor
      1 bubblorna
      1 bubblornas
      1 bubers
      1 buboner
      2 bubonerna
      1 bud
      4 budbärare
      1 buddchiari
      1 buddha
      1 buddhism
      6 buddhismen
      2 buddhismens
      1 buddhisten
      1 buddhistisk
      5 buddhistiska
      1 buddhistiskthinduistiska
      1 buddhistmunkar
      1 buddismen
      1 budgeten
      1 budgetklass
      1 budo
      1 budouövare
      1 buds
      1 budskap
      1 budskapet
      1 buffalo
      1 buffer
      4 buffertens
      4 buffertformeln
      1 buffertlösning
      1 buffertsystem
      1 buffertverkan
      1 buffra
      1 buffrande
      1 buffras
      1 buffycoat
      2 bugchasing
     10 buk
      1 bukandningen
      1 bukaorta
      1 bukaortaaneurym
      5 bukaortaaneurysm
      1 bukarest
      1 bukarna
      1 bukduk
     53 buken
      1 bukens
      1 bukfenorna
     34 bukfetma
      2 bukfetman
      3 bukhåla
     21 bukhålan
      8 bukhinnan
      1 bukhinnedialys
      1 bukhinnehålan
      6 bukhinneinflammation
      1 bukhinneinflammationen
      1 bukhinneöverdrag
      1 bukhinnevävnad
      1 bukhuden
      2 bukinfektioner
      1 bukinnehållet
      1 bukkirurgin
      1 bukmuskler
      1 bukmusklerna
      3 bukmuskulaturen
      1 bukområdet
      2 bukoperation
      1 bukoperationerna
      1 bukorganen
      4 bukplastik
      2 bukplastiken
      1 bukröntgen
     10 buksmärta
      1 buksmärtan
      9 buksmärtor
      2 buksnitt
      4 bukspott
      1 bukspottet
      5 bukspottkörtel
      1 bukspottkörtelcancer
      7 bukspottkörtelinflammation
     25 bukspottkörteln
      3 bukspottkörtelns
      1 bukspottskörtelgången
     11 bukspottskörteln
      2 bukspottskörtelns
      1 bukspottskörtlar
      1 bukspöttskörtlar
      5 bukt
      1 bukta
      4 buktar
      1 bukter
      1 buktryck
      1 bukvägg
     16 bukväggen
      1 bula
      2 bulak
      1 bulber
      1 bulbiller
      1 bulbocodium
      2 bulgarien
      1 bulges
      1 bulimi
      5 bulimia
      2 buljong
      4 bulkmedel
      3 bull
      1 bullan
     27 buller
      1 bullerdämpning
      1 bullerexponeringen
      1 bullerkällan
      1 bullermätning
      3 bullernivå
      2 bullerplank
      1 bullerreducerande
      1 bullerreducering
      1 bullersänkande
      1 bullerskadade
      3 bullerskador
      1 bullerutsläckning
      1 bullerutsläppen
      1 bulleryrkena
      1 bulletin
      1 bullionmynt
      2 bullös
      1 bullrande
      4 bullret
      3 bullriga
      1 bullsfoot
      3 bulor
      1 bultning
      1 bumps
     15 bunden
      1 bundenhet
      2 bundesamt
     15 bundet
      1 bundibugyo
      1 bundistammen
      6 bundit
      4 bundna
      1 bunke
      1 bunt
      2 buntar
      1 bunyan
      1 bunyavirus
      1 bup
      1 buprenorfin
      1 burbridge
      2 burden
      3 buren
      4 burgdorferi
      1 burghardt
      2 burit
      2 burk
      1 burka
      1 burkar
      1 burkholderia
      1 burkitts
      1 burma
      1 burned
      1 burnet
      1 burnetii
      6 burnetti
      1 burows
      3 bursa
      2 bursit
      1 burton
      2 burundi
     12 buskar
      1 buskarna
      6 buske
      1 buskens
      1 buskig
      1 buskilla
      1 buskliknande
      1 buskmarker
      1 busnh
      1 busnsnbu
      4 buss
      1 bussanalysator
      1 bussarong
      2 bussen
      1 bussspårvagnsförare
      1 bussy
      1 büstenhalter
      1 busters
      1 bustiern
      1 bustiers
      1 butenandt
      1 butik
      1 butiken
      7 butiker
      2 butler
      1 butylgruppen
      1 butylhydroxianisol
      1 butylkedjor
      1 butyrospermum
      2 bv
      1 bviruskodat
      1 bvitaminbesläktade
      4 bvitaminer
      1 bvitaminerna
      1 bvitaminet
      1 bvitaminkomplexet
      6 by
      5 byar
      1 bybor
      1 byfånarna
      2 bygdemål
      1 bygdens
      5 bygel
      1 bygelbehåar
      2 bygelbh
      1 bygeln
      1 bygg
     19 bygga
      1 byggämnesmaterial
      1 byggande
      2 byggandet
      1 byggarbetssamordnare
      7 byggas
      1 byggbranschen
      2 byggd
      1 byggda
      7 byggde
      5 byggdes
     68 bygger
      1 byggindustrin
      1 bygglagen
      1 bygglov
      1 byggmaterial
      9 byggnad
      2 byggnaden
     11 byggnader
      1 byggnadsägaren
      1 byggnadsakustik
      1 byggnadsämnesindustri
      1 byggnadsarbetare
      2 byggnadskonst
      3 byggnadsmaterial
      1 byggnadsminnesmärkt
      1 byggnadssätt
      1 byggnadsställning
     14 byggs
      4 byggsten
      6 byggstenar
      6 byggt
      6 byggts
      1 byggvaruhus
      2 byglar
      1 byglarna
      1 byk
      1 byläkare
      1 byling
      4 byn
      1 byns
      2 bypass
      1 bypasskirurgi
      1 byprästen
      2 byråkratiska
      2 bysantinska
      8 byst
      1 bystdrottningarna
     21 bysten
      2 bysthållare
      1 bystomfånget
      2 byt
     29 byta
     12 bytas
     20 byte
     12 byten
      1 bytena
      8 byter
      5 bytesdjur
      3 bytesdjuret
      1 bytesdjurets
      6 bytet
     19 byts
      5 bytt
     11 bytte
      4 byttes
      1 bytts
      1 byxfickan
      1 byxgalge
      1 byxmyndighetsåldern
      3 byxor
     78 c
     62 �c
      6 ��c
    181 ca
      1 cabrerianus
      1 cachexia
      2 cacl
      1 caclclo
      1 cacl[clo]
      2 caclo
      2 caco
      1 cadherincateninkomplex
      1 cadmium
      1 cadolle
      1 cadolles
      3 caecum
      1 caedare
      2 caesar
      1 caesarea
      1 caesars
      1 caeso
      1 caféaulaitfärgad
      1 caféaulaitfläckar
      1 caffeinated
      1 caffeine
      1 cag
      3 cage
      1 cahco
      1 cairns
      1 caivano
      1 cajal
      1 cajalretziusneuroner
      1 cakra
      1 calais
      2 calcgenen
      1 calculus
      1 calea
      1 calibur
      6 calicivirus
      2 california
      2 californicum
      1 callahan
      1 callosotomi
      1 calls
      2 calmette
      2 calmetteguérin
      1 calor
      1 caloric
      1 calorie
      2 calycibus
      1 cam
      6 cambridge
      1 cambridgekuren
      2 cambridgemåltider
      1 cambrige
      1 camgfesiooh
      2 camille
      1 camillo
      1 campbell
      1 campestris
      1 camping
      1 campingplatser
      1 campos
      1 campus
      4 campylobacter
      1 camus
      1 can
      4 canada
      2 canadensis
      1 canadian
      1 canalis
      1 canberra
    234 cancer
      6 cancerbehandling
      4 cancercell
      3 cancercellen
     22 cancerceller
      2 cancercellerna
      2 cancercellstypen
      1 cancerdiagnos
      1 cancerdödsfallen
      1 cancerdrabbad
      5 cancerfall
      1 cancerfallen
      2 cancerfonden
      4 cancerform
      8 cancerformen
     18 cancerformer
      1 cancerformerna
      1 cancerforskningen
      1 cancerforskningsinstitut
      1 cancerframkallade
     14 cancerframkallande
      1 cancergener
      1 cancerhämmande
      1 cancerhundar
      1 cancerinsjuknanden
      1 cancerknölar
      1 cancerläkaren
      1 cancerliknande
      2 cancermarkör
     29 cancern
      1 cancerns
      3 cancerogen
      1 cancerogena
      3 cancerogent
      1 cancerorksaken
      1 cancerösa
      1 cancerpatient
      1 cancerpatienten
      4 cancerpatienter
      1 cancerrelaterade
      3 cancerrisk
      1 cancerrisken
      1 cancersjuk
      6 cancersjukdom
      5 cancersjukdomar
      1 cancerspridning
      1 cancerstadiet
      1 cancerstamceller
      1 cancersvulster
      1 cancerterapi
      1 cancertumören
      3 cancertumörer
      3 cancertyp
      2 cancertypen
      3 cancertyper
      2 cancerunionen
      1 canceruppkomst
      1 cancerupptäckt
      1 cancerutredning
      1 cancerutveckling
      1 cancervård
      1 cancervävnad
      7 cancrar
      8 candida
      1 candide
      3 candidiasis
      1 candidosis
      1 canetti
      1 canine
      1 canines
      2 canis
      1 cannabiod
     36 cannabis
      2 cannabisanvändning
      2 cannabisbruk
      1 cannabisbruket
      1 cannabisbrukets
      1 cannabiscigaretter
      1 cannabisfolket
      4 cannabisrökning
      1 cannes
      1 cannies
      1 cannula
      1 cant
      1 cantonensis
      2 cantor
      1 cao
      1 caoh
      1 cap
      1 capablanca
      1 capacitet
      2 capacity
      1 capgras
      2 capitis
      1 caplan
      2 capooh
      1 capsaicintest
      2 capsulatum
      1 caput
      1 cara
      1 caramanicum
      3 carateum
      1 caravaggio
      2 carb
      1 carcinoembryogent
      1 carcinogen
      1 carcinogena
      3 carcinogener
      1 carcinogenes
      1 carcinoid
      1 carcinoida
      1 carcinoidsyndrom
     41 carcinom
      4 carcinoma
      1 carcinomatofobi
      1 carcinomatos
      2 carcinomet
      1 carcinomgruppen
      1 cardia
      1 cardiale
      1 cardinalhealth
      1 cardiolite
      1 cardiovascular
      3 care
      1 carin
      2 carinatum
      1 carinatus
      1 cariniiinfektioner
     20 carl
      1 carla
      2 carlbeck
      1 carlgustav
      1 carlo
      1 carloscar
      1 carlsen
      7 carlsson
      1 carlström
      1 carmichaelii
      1 carney
      1 carniolica
      1 carnivore
      1 carnivorer
      1 carol
      3 carolina
      1 caroline
      2 caroticus
      1 carpaccio
      1 cars
      1 carseywerner
      1 cartilagines
      4 cartilago
      2 carukia
      1 caruncula
      1 casciarolus
      1 casebook
      2 casecontrol
      1 casereferent
      1 casey
      1 cashew
      1 cashewnötter
      1 casnr
      2 casnummer
      1 caso
      1 caspar
      1 caspofungin
      2 cassette
      1 cassidy
      1 cassius
      1 castaway
      1 castrare
      1 castren
      1 casts
      7 cat
      1 catalepsis
      7 catalogue
      2 catarina
      2 catarrhalis
      1 catathrenia
      4 catch
      4 catgut
      1 catgutet
      1 catguts
      2 catguttrådarna
      1 catharanthus
      1 catharina
      1 catherine
      1 cathéter
      1 cativaprocessen
      1 cattell
      1 cattells
      1 cattellskalan
      1 cauchemar
      1 cauda
      1 caudatum
      1 causis
      1 cauv
      5 cava
      1 cave
      1 cavernosa
      1 cavum
      1 cayennepeppar
      2 cb
      2 cbct
      1 cbd
      1 cbs
      1 cce
      1 cceller
      2 ccellerna
      1 ccim
      5 cck
      1 cckpeptiden
      1 cckpeptider
      1 cckpz
      1 ccks
      3 ccu
     11 cd
      4 cdc
      1 cdcellerna
      1 cdco
      1 cdh
      1 cdmolekyl
      1 cdmolekylen
      1 cdna
      1 cdproteiner
      1 cdrom
      2 cds
      1 cdspecifik
      1 cdspelare
      1 cdsupermab
      2 cdtal
      2 cdtekniken
      2 ce
      2 cea
      1 cecum
      1 cederträd
      2 cefalexin
      1 cefalgi
      2 cefalosporin
      1 cefalosporinantibiotika
     13 cefalosporiner
      1 cefalosporinpreparat
      2 cefic
      2 cefotaxim
      6 ceftriaxon
      1 celebra
      2 celebriteter
      4 celecoxib
      1 celgene
      1 celiaker
     26 celiaki
      1 celibat
     25 cell
      4 celladhesion
      1 celladhesionen
      1 celladhesionsmolekyler
      1 cellager
      1 cellandning
      3 cellandningen
      3 cellanemi
      1 cellantalet
      1 cellbundna
      1 cellcykelhämmare
      2 cellcykeln
      1 cellcykelns
      1 celldelas
     23 celldelning
      4 celldelningar
      2 celldelningarna
      1 celldelningen
      1 celldifferentiering
     15 celldöd
     61 cellen
      1 cellenreceptorn
     15 cellens
    248 celler
      2 �celler
      1 cellerdygn
      1 cellerl
     73 cellerna
      8 cellernas
      1 cellerul
      1 cellförändring
      1 cellförändringar
      1 cellförbindelserna
      2 cellform
      1 cellformer
      1 cellforskaren
      1 cellfragment
      8 cellgift
     16 cellgifter
      1 cellgifts
      1 cellgiftsbehandlig
      8 cellgiftsbehandling
      1 cellgiftsbehandlingen
      1 cellhämmande
      1 cellhämmare
      1 cellini
      1 cellinnehåll
     11 cellkärna
      2 cellkärnan
      2 cellkärnor
      1 cellkärnornas
      1 cellklump
      7 cellkroppen
      1 celllära
      1 cellmassa
      1 cellmassan
      1 cellmaterial
      1 cellmedierad
     18 cellmembran
      2 cellmembraner
     22 cellmembranet
      1 cellmembranfunktion
      1 cellmetabolismen
      1 cellmodeller
      1 cellnedbrytning
      1 cellnekros
      4 cellnivå
      1 cellnybildning
      2 cellodling
      2 cellodlingar
      2 cellomsättning
      2 cellplasma
      3 cellplasman
      1 cellpopulationen
      1 cellproduktion
      1 cellproliferation
      2 cellprov
      1 cellprover
      1 cellreproduktionen
      2 cells
      2 cellskräck
      1 cellsträng
      1 cellstruktur
      1 cellterapier
      5 celltillväxt
      1 celltillväxthämmande
      1 celltoxiskt
      5 celltyp
      1 celltypen
      5 celltyper
      1 celltyperna
      1 cellular
      3 cellulär
      2 cellulära
      1 cellularpathologie
      2 cellulärt
      1 cellulin
      5 cellulit
      1 cellulite
     11 celluliter
      3 celluliterna
      1 cellulitis
      1 celluloidplåtar
      6 cellulosa
      1 cellulosaacetat
      1 cellulosaacetatbågar
      1 cellulosafibrerna
      2 cellulosamaterial
      1 cellulosan
      1 cellulosanitrat
      1 cellulosapropionat
      2 cellulosapropionatbågar
      1 cellulosapulver
      1 cellutbyte
     16 cellvägg
      1 cellväggar
      7 cellväggen
      1 cellvandring
      1 cellvävnad
      1 cellvävnader
      1 cellvibrationer
      6 cellytan
      3 cellytor
     13 celsius
      6 celsus
      2 cemärkning
      5 cement
      1 cementen
      1 cementsealer
      1 cengage
      1 centc
      4 center
      7 centers
      1 centesimalpotensen
     68 centimeter
      7 centimeters
      1 centimeterstora
      1 centimeterstorlek
      5 centra
      1 centrakstimulerande
     45 central
    151 centrala
      2 centralafrika
      4 centralafrikanska
      4 centralamerika
      4 centralasien
      1 centralbanker
      2 centralbyrån
      4 centraleuropa
      1 centralförbundet
      1 centraliserad
      1 centralisering
      1 centrallasarett
      1 centralsjukhus
      3 centralstimulantia
      1 centralstimulerade
     11 centralstimulerande
     18 centralt
      3 centre
      2 centrerad
      1 centrerade
      1 centret
      1 centrifuger
      1 centrifugera
      1 centrifugerar
      1 centrifugeras
      1 centrosom
     25 centrum
      1 centrumet
      1 centrumfrekvensen
      1 centurioner
      2 cephenemyia
      2 cerat
      1 cerea
      2 cerebellum
     13 cerebral
      3 cerebrala
      1 cerebralt
      1 cerebri
      1 cerebrospinal
      1 cerebrospinalis
     12 cerebrospinalvätska
     13 cerebrospinalvätskan
      1 cerebrovaskulära
      1 ceremoniella
      2 ceremonier
      1 ceremonin
      3 cereus
      1 cerkariedermatit
      1 cerkarier
      2 cerkarierna
      1 cerkarium
      1 cerremonikaraktär
      1 certifiera
      3 certifierade
      2 certifierat
      2 certifiering
      1 certifieringsprov
      1 certifikat
      8 ceruloplasmin
      1 ceruloplasminprotein
      1 cervarix
      1 cervi
      1 cervical
      2 cervicit
      1 cervikal
      2 cervix
      4 cervixcancer
      1 cervixpessar
      1 cesarea
      3 cescau
      2 cesium
      2 ceskoslovensk�
      1 cetera
      1 cetylpyridin
      6 cetylpyridinklorid
      2 cf
      1 cfc
      1 cformad
      3 cfuml
      1 cgm
     17 ch
      1 chagas
      3 chain
      1 chairman
      6 chakra
      1 chakrabalansering
      1 chakraläran
      6 chakran
      1 chakras
      2 chakrasystemet
      1 chakror
      1 chamber
      1 chamberland
      1 chamberlen
      1 chamboning
      1 champagneflaska
      1 champna
      1 champo
      1 chanel
     18 chans
      5 chansen
      4 chanser
      7 chanserna
      2 chapel
      1 characteribus
      2 characteristics
      1 characterization
      1 charak
      1 charaka
      2 charakas
      1 charge
      1 charifloden
      2 charité
      1 chark
      2 charken
      2 charker
      1 charlatan
      1 charlatanen
     16 charles
      2 charlesbogerti
      1 charlotta
      3 charlotte
      4 charm
      2 charmen
      1 charmerande
      1 charmören
      2 charri�re
      2 chasing
      5 chastel
      1 chastels
      1 chato
      1 chatta
      1 chattar
      1 chauliac
      2 chazes
      3 chbr
      1 chchchoh
      1 chchnh
      2 chchoh
      5 chcl
      1 chclcooh
      2 chclf
      1 chcln
      2 chclnop
      1 chclnos
      3 chclo
      1 [chco]o
      3 chcooh
      1 checkboxar
      1 checklista
      1 checklistan
      2 checklistor
      6 chef
      5 chefer
      1 chefredaktör
      1 chefstjänsteman
      1 chefstjänstemannen
      1 cheir
      1 chek
      1 chelidonium
      5 chemical
      2 chemicals
      1 cheney
      2 cheopis
      1 cher
      1 cherry
      1 chesebroughponds
      1 chester
      1 chewing
      1 chfnos
      4 chi
      2 chiapas
      1 chicago
      4 chief
      1 chihuahua
      3 chikungunya
      1 child
      3 children
      4 chile
      1 chilesalpeter
      1 chillums
      2 china
      1 ching
      1 chiro
      1 chironex
      3 chiropractic
      1 chiropraktorsällskapet
      1 chiti
      1 ch�jio
      8 chlamydia
      5 chlamydophila
      1 chloromycetin
      3 chls
      4 chn
      2 chncl
      1 chnh
     10 chno
      6 cho
     36 chock
      1 chockartad
      1 chockterapi
      1 chocktillstånd
      1 chockvågor
      2 chockvågsbehandling
     13 choh
      1 chohcooh
      1 choho
     10 choklad
      1 chokladen
      4 chokladförgiftning
      1 chokladprodukter
      1 cholangiocarcinom
      1 cholangiocarcinoma
      5 cholecystektomi
      5 cholecystit
      1 cholecystokinin
      1 choledochi
      4 choledochus
      1 cholerae
      1 cholestasislymphedema
      1 cholesystokinin
      2 cholsyra
      1 chon
      1 chona
      1 chondrus
      1 chongzhen
      1 chooh
      1 chorda
      5 chorea
      1 chorioretinalt
      1 chorioretinit
      1 choroidea
      3 choroideus
      1 chos
      1 chovsteks
      1 chrétien
      1 chris
      1 christer
      1 christiaan
      9 christian
      1 christmas
      7 christopher
      1 chroma
      1 chromolaena
      1 chronic
      1 chronically
      1 chronicle
      1 chronicum
      1 chronicus
      1 chrysanthus
      1 chrysogenum
      1 chsn
      1 chso
      1 chungs
      1 church
      1 chürgstrauss
     11 chymus
      3 ci
      3 cia
      1 cialis
      1 ciao
      1 cicuta
      1 cider
      5 cigarett
      1 cigarettdimma
      6 cigaretten
     15 cigaretter
      2 cigarettes
      1 cigarettetuier
      1 cigarettfilter
      1 cigarettmarknaden
      1 cigarettmunstycken
      8 cigarettrök
      3 cigarettrökning
      1 cigarr
      2 cigarren
      7 cigarrer
      1 cigarrlåda
      1 cigarrlådor
      1 cigarrsnoppare
      1 cihuacoahuatl
      1 ciimplantat
      1 cikador
      2 ciliare
      1 ciliarmuskeln
      1 ciliarmuskelspänningen
      1 ciliarnerverna
      1 cilicicus
      1 cilie
      2 cilier
      1 cilierade
      3 cilierna
      1 ciliolatus
      7 cimex
      1 cinctum
      1 cinerea
      1 cingulate
      1 cinguli
      1 cingulin
      1 cinhibitor
      1 cinhibitorkoncentrat
      1 cinnober
      1 ciofis
      1 cioms
      1 ciopereras
      1 cip
      1 cipav
      1 cipro
      5 ciprofloxacin
      1 ciproxin
      1 circuit
      1 circumforaneos
      2 circumventrikulära
    337 cirka
      3 cirkel
      1 cirkelbåge
      1 cirkelrund
      1 cirkelrunda
      1 cirkelträning
      3 cirkulära
      1 cirkulärt
      6 cirkulation
      9 cirkulationen
      2 cirkulations
      1 cirkulationseffekt
      1 cirkulationshämmande
      1 cirkulationsinsufficiens
      2 cirkulationskollaps
      1 cirkulationsluft
      1 cirkulationsorganen
      2 cirkulationsplats
      2 cirkulationsrubbningar
      1 cirkulationsstillestånd
      1 cirkulationsstimulerande
      7 cirkulationssvikt
      1 cirkulationssymtom
      2 cirkulationssystem
      4 cirkulationssystemet
      2 cirkulatorisk
      2 cirkulatoriska
      2 cirkulera
      8 cirkulerande
     12 cirkulerar
      2 cirkumpolär
      1 cirkus
      1 cirrhosis
      1 cirrhosus
      3 cirros
      2 cirrosens
      1 cis
      1 citalopram
      2 citat
      1 citaten
      1 citerats
      3 cites
      2 citodon
      4 citrat
      2 citron
      1 citronellol
      1 citronsaft
      5 citronsyra
      4 citronsyracykeln
      1 citrusfrukt
      2 citrusfrukter
      3 city
      6 civil
     12 civila
      1 civilbilar
      1 civilisationen
      4 civilisationer
      1 civilisationerna
      1 civilklädda
      1 civilplikt
      1 civilrätt
      3 civilrättslig
      4 civilrättsliga
      1 civilstånd
      1 civilt
      1 cj
      1 ckit
      1 cknivån
      1 ckupa
      1 cl
      1 cla
      1 cladosporium
      1 claes
      1 claforan
      1 claq
      1 claritromycin
      1 clarity
      1 clark
      1 class
      1 classical
      5 classification
      1 claude
      2 claudicatio
      1 claudiner
      1 claudio
      1 claustrophobia
      1 claustrum
      3 claviceps
      9 clearance
      1 clearancen
      1 clearancer
      1 clearancerna
      3 clearleft
     42 clearright
      3 cleckley
      1 cleland
      1 clematitis
      1 clemens
      1 clermontferrand
      1 clethra
      1 cliffs
      1 clinic
      4 clinical
      1 clinicla
      2 clinique
      2 clips
      1 clitoris
      1 clitorism
      1 cll
      1 clo
      1 clofazimin
      1 clonal
      1 closener
      1 closeness
     11 clostridium
      1 clostridiumarter
      1 clover
      1 club
      1 cluny
      1 clutter
      1 cluttons
      1 clv
      1 clymenum
      1 clynes
     95 cm
      6 �cm
      1 cm�
      1 cmax
      1 cmbred
      2 cmho
      2 cmv
      1 cmvinfektion
      2 cn
      1 cn�
      1 cnd
      1 cnhnmohm
      1 cnhon
      1 cnidaria
      1 cnidocyt
      1 cnidocytes
      1 cnnh
      6 cns
     14 co
      2 coacher
      1 coagonist
      1 coahuila
      2 coast
      1 cobain
      3 cobb
      2 coca
      1 cocacola
      2 coccidioides
      1 coccidioidomykos
      5 cochleaimplantat
      2 cochlean
      6 cochrane
      1 cochranes
      1 cocillana
      1 cocktailar
      1 coding
      1 codrington
      1 coenzym
      2 coeruleus
      4 coeundi
      1 coffee
      1 cogmed
      3 cognitive
      1 cohalten
      1 cohen
      1 coherence
      1 cohesivgelproteser
      1 cohors
      1 cohortes
      1 coinfektion
      1 coitus
      2 cola
      1 colchicin
      1 colchicinet
      3 colchicum
      1 colchicumarterna
      2 cold
      1 coldplay
      1 coleman
      3 colgate
      4 colgatepalmolive
     16 coli
      1 colin
      1 colit
      2 collaboration
      3 college
      1 collegiet
      6 collegium
      1 colliculus
      1 collie
      1 collip
      3 colombia
      1 colombiansk
      7 colon
      1 coloningjutning
      1 colonkolon
      2 colorado
      1 colostomi
      1 coltsfoot
      1 columbian
      1 columbianhypotesen
      2 columbinemassakern
      1 columbit
      1 columbus
      1 columbusresa
      1 colworth
      1 com
      5 coma
      2 comar
      1 comättnaden
      2 come
      4 comfort
      1 comics
      1 comité
      1 commercial
      4 commission
      1 commitment
      4 committee
      1 committeé
      1 committment
      4 common
      2 commotio
      2 communication
      2 communications
      3 communis
      1 communisse
      3 community
      1 comorbidity
      2 compact
      6 company
      1 compartmentsyndrom
      1 complete
      2 complex
      3 compliance
      1 compound
      1 comprehensive
      1 compulse
      1 computational
      2 computed
      1 computers
      1 comt
      1 con
      1 concept
      1 concerta
      1 conditionett
      1 conditions
      1 conduct
      1 condyline
      2 condyloma
      1 conference
      1 congar
      1 congelatio
      1 congenita
      1 congenital
      1 congolese
      1 conh
      1 conicae
      1 conidae
      1 conjugated
      3 connecticut
      1 connelly
      1 conneticut
      1 connors
      3 conns
      1 conoclinium
      1 conotruncal
      1 conquistadorerna
      1 conrad
      1 consciousness
      1 conservative
      1 considerable
      8 consortium
      1 consortiums
      1 constabulary
      1 construction
      1 consumer
      1 consumers
      1 contagiosa
      1 containerdykning
      1 containrar
      1 contergan
      5 continuous
      4 contorix
      1 contortatall
      2 contortrix
      1 contre
     13 control
      1 controlled
      1 controlprogrammet
      1 convallaria
      1 convallariaceae
      1 convallium
      1 convention
      1 converting
      1 convulsive
      1 conyzoides
      2 cooke
      1 cooköarna
      1 cooks
      2 coombs
      1 cooper
      1 coordination
      1 coover
      1 copco
      1 copd
      3 cope
      2 coping
      2 copingstrategi
      2 copingstrategier
      1 copp
      1 copulatio
      1 copulerades
      1 copulerakopulera
      8 copycat
      1 copycatbrott
      1 copycatbrotten
      2 copycatbrottet
      1 copycatbrottslingar
      1 copycateffekt
      2 copycateffekten
      1 copycaten
      1 copycats
      1 copying
      1 cord
      1 cordis
      1 core
      3 coricykeln
      2 corioliseffekten
      1 cornea
      2 cornell
      1 corneum
      2 cornutum
      5 corona
      4 coronavirus
      1 coronaviruset
      1 corpora
      1 corporation
      2 corporis
      1 corpulence
     14 corpus
      1 correlation
      1 cors
      1 corset
     11 cortex
      3 cortiska
      1 corvisart
      1 corylifolia
      1 corynebacterium
      3 cosby
      1 cost
      1 costales
      1 couldnt
      9 council
      2 couney
      1 counseling
      2 counterblaste
      1 countries
      2 county
      1 couple
      1 courage
      1 court
      1 courtois
      1 cousin
      3 couvade
      2 couver
      1 couveuse
      1 covidien
      1 cowboyen
      1 cowpers
      3 cox
      3 coxiberna
      3 coxiella
      1 coyette
      1 cp
     22 cpap
      2 cpapanvändare
      2 cpapapparat
      2 cpapapparaten
      2 cpapapparater
      1 cpapbehandling
      1 cpapmaskin
      1 cpatienter
      2 cpeptid
      1 cpeptiden
      3 cpg
      1 cpim
      1 cpk
      1 cpotenser
      2 cpskada
      3 crack
      1 craps
      1 crash
      1 craske
      2 crassum
      1 craving
      1 crawford
      1 creaktioner
      1 creaktiv
      4 creaktivt
      1 credé
      1 credés
      1 credit
      1 credits
      1 cremaster
      2 cremastermuskeln
      1 creme
      1 cremefärgade
      1 cremeliknande
      1 cremello
      1 crescentnefrit
      1 crestor
      1 crétin
      3 creutzfeldtjakobs
      2 creutzfeldt�jakobs
      1 cribrosa
      1 crichton
      1 crick
      1 cricket
      1 cricoarytenoidmuskeln
      1 cricofaryngeus
      2 cricoidea
      1 crispus
      2 critical
      1 critonia
      2 cro
      1 crocparytenoidmuskeln
      1 croft
      1 croghan
      1 crohn
      8 crohns
      1 crosby
      1 crosscut
      1 crotalus
      1 crow
      8 crp
      1 crptest
      1 crt
      1 cru
      1 crüe
      1 cruise
      2 cruris
      1 crus
      1 crusta
      1 cruzi
      1 cryonics
      2 cryonite
      1 cryoniten
      2 cryptococcus
     24 cryptosporidium
      1 cryptosporidum
      1 cryptostegia
      1 crystallized
      2 csf
      1 csns
      3 css
     20 csv
      1 csvanalysen
      1 csvflöde
      1 csvglukos
      1 csvglukosvärdet
      1 csvläckage
      1 csvodlingen
      1 csvprovet
      1 csvvärdena
      9 ct
      1 ctbilder
      1 ctcomputer
      1 c�te
      1 ctg
      1 cttft
      1 cubare
      1 cubomedusae
      1 cubozoa
      1 cuitlacochi
      2 culex
      1 culicidae
      2 culicinae
      1 culiseta
      1 cullen
      1 cultural
      2 cum
      1 cumbia
      1 cummingtonit
      1 cunninghams
      1 cupping
      2 cura
      1 curaisserespiratorer
      1 curare
      1 curbpoängen
      2 curcumin
      1 curcuminoiden
      1 curcuminoiderna
      4 curentur
      3 curie
      1 curieinstitutet
      1 curies
      1 curman
      2 curt
      2 curvatura
      2 curve
      1 cuscuta
      1 cushing
     10 cushings
      3 cuspen
      1 cutis
      1 cutting
      1 cuvilliers
      1 cuzco
      1 cvapenarsenaler
      2 cvd
      1 cvddiagnosen
      8 cvitamin
      1 cvitaminbrist
      1 cvitaminets
      1 cvitaminpreparaten
      1 cvitaminrik
      1 cvk
      1 cvl
      1 cvsymmetri
      1 cvz
      1 cyan
      1 cyanamid
      1 cyaneus
      1 cyanhaltiga
      6 cyanid
      1 cyanidalstrande
      2 cyanider
      1 cyanidförgiftning
      1 cyanidjonen
      2 cyanoacrylat
      1 cyanoacrylatlim
      1 cyanoakrylat
      1 cyanoakrylsyra
      1 cyanogen
      1 cyanogeniska
      1 cyanopropensyra
     19 cyanos
      1 cyanotisk
      1 cyansyra
      1 cyanväte
      1 cyanväteförgiftning
      1 cybernetisk
      2 cyborg
      4 cyborger
      1 cyclodehydration
     11 cykel
      1 cykelbana
      2 cykelbanor
      1 cykelbyxor
      1 cykelfält
      1 cykelhandbromshandtag
      8 cykeln
      1 cykelpedaler
      1 cykelrunda
      1 cykelväg
      1 cykla
      2 cyklar
      4 cykler
      1 cyklerna
      2 cykling
      4 cyklisk
      4 cykliska
      4 cykliskt
      1 cyklist
      1 cyklisten
      3 cyklister
      1 cykloadditionen
      1 cykloalkaner
      7 cyklofosfamid
      1 cyklohexan
      3 cyklohexanol
      4 cyklohexanon
      2 cyklohexanring
      2 cykloheximid
      2 cykloid
      1 cyklokapron
      1 cyklonit
      1 cyklooxgenas
      1 cyklopropen
      1 cyklotron
      4 cyklotymi
      1 cyklotymier
      1 cyl
      2 cylinder
      1 cylinderceller
      3 cylinderepitel
      1 cylinderepitelet
      1 cylinderformade
      1 cylinderglas
      1 cylindern
      3 cylindrisk
      5 cylindriska
      2 cylindriskt
      1 cynapium
      1 cynisk
      2 cyp
      2 cypa
      1 cypc
      5 cypern
      2 cypgener
      1 cyritestin
      1 cyst
     13 cysta
      5 cystan
      1 cystans
      1 cystatin
      1 cystbildning
      1 cysteinrikt
      1 cysteinylleukotrien
      1 cystform
      1 cystformen
      2 cystica
      1 cysticercos
      1 cysticerkos
      4 cysticus
      2 cystinsten
      1 cystinstenar
     11 cystisk
      2 cystiska
      1 cystiskt
      4 cystit
      1 cystitis
     19 cystor
      1 cystorkan
      2 cystorna
      1 cystornas
      2 cystoskop
      3 cystoskopi
      1 cystostaticum
      2 cytalidium
      1 cytarabin
      1 cytisin
      1 cytogena
      1 cytogenetisk
      2 cytokin
     20 cytokiner
      1 cytokinet
      1 cytokininducerad
      1 cytokininer
      2 cytokrom
      3 cytologi
      1 cytologisk
      3 cytologiska
      4 cytomegalovirus
      1 cytomegalovirusretinit
      8 cytoplasma
      1 cytoplasmaenzymer
      5 cytoplasman
      1 cytoplasmiska
      1 cytoskelettet
      1 cytoskopi
      1 cytosol
      2 cytosolen
     28 cytostatika
      3 cytostatikabehandling
      2 cytostatikum
      1 cytotoxisk
      1 cytotoxiskt
      1 czeczottianus
     58 d
     11 da
   1564 då
      1 dä
      1 daao
      1 daboia
      1 dachau
      1 däck
      6 dadamo
      1 dadamos
      1 dafrisättningen
    166 dag
      2 daga
    197 dagar
      1 �dagar
     18 dagarna
      1 dagarref
      9 dagars
      1 dagdrömmer
     55 dagen
     61 dagens
      1 daggblå
     76 däggdjur
      3 däggdjuren
      4 däggdjurens
      2 däggdjurs
      2 däggdjursarter
      1 däggdjurshonor
      1 däggdjursinsulin
      1 däggdjursordningar
      4 daggmaskar
      1 daggmaskarnas
      1 daggmaskens
      1 daghem
      1 dagis
      1 dagisvistelse
      8 daglig
     24 dagliga
     21 dagligen
     32 dagligt
      2 dagligvaror
      1 dagligvaruaffärer
      1 dagligvarubutiker
      3 dagligvaruhandel
      1 dagligvaruhandeln
      1 dagnos
      1 dagordning
      8 dags
      1 dagsböter
      9 dagsläget
      1 dagsljus
      1 dagsljuslysrör
      1 dagstidningar
      1 dagsymptomen
      9 dagtid
      1 dagtidssymptom
      2 dagtrötthet
      1 dagtröttheten
      1 daguerrotypi
      1 dagvis
      1 dahlberg
      1 dahlin
      1 dahlstedt
      2 daigremontianum
      2 dairy
      7 daisy
      3 daisyböcker
      1 daisybok
      2 daisyformatet
      1 daisyformatets
      1 daisyprogramvara
      1 daisyspecifikation
      1 daisyspecifikationer
      3 daisyspelare
      1 daktulos
      1 daktylisk
      1 dala
      1 dalälven
      1 dalälvens
      4 dalanin
      5 dalaninrest
      1 dalaninresten
      1 dalaninstrukturen
      5 dalarna
      1 dale
      1 dalgång
      1 dalgångar
     90 dålig
     20 dåliga
     56 dåligt
      1 dallas
      1 dallilja
      1 dallrar
      3 dalsland
      3 dalton
      1 dam
      1 damascena
      1 damaskus
      1 dambågar
      1 dambinda
      1 dame
      1 damer
      1 damerna
      1 damers
      1 damfetaminsalt
     11 damm
      3 dammar
      1 dammet
      1 dammfria
      5 dammlunga
      1 dammpartiklar
      3 dammsuga
      2 dammsugare
      2 dammsugaren
      1 dammsugning
      1 dammtorkning
      1 damocratis
      2 damokrates
     14 damp
     16 dämpa
      1 dämpad
      1 dämpade
      1 dampadhddiagnostiken
      9 dämpar
      3 dämpas
      1 dämpning
      1 dämpningen
      1 damsugare
      1 damulstertyg
      1 damunderkläder
      1 damunderplagg
      1 dan
      1 dana
      1 danas
      2 danazol
      1 danderyds
      3 dandy
      1 dandyfeber
      2 danert
      3 daniel
      2 dänkflaskor
      2 danlos
     37 danmark
      1 danmarks
      1 danocrine
      4 dans
      2 dansa
      1 dansade
      1 dansande
      2 dansare
      1 dansarna
      1 dansbaserad
      1 dansbaserade
      2 dansen
      1 danser
      2 danshantlar
      1 dansimpuls
      3 dansk
      4 danska
      1 danskan
      1 danskans
      3 danske
      1 danskonsten
      1 danskoreografi
      2 danskt
      1 danslärare
      1 dansmani
      3 danssjuka
      1 danssjukan
      1 danssko
      1 danssneaker
      1 danssteg
      1 dao
      4 daphne
      1 daphnetoxin
      2 dapson
      1 daptomycin
   1316 där
     40 därav
    154 därefter
      2 däremellan
    155 däremot
    527 därför
      6 däri
     52 däribland
     24 därifrån
     61 därigenom
      1 därinne
      2 därjämte
      1 dark
      1 darkness
      1 darling
    238 därmed
      2 därom
      4 dårört
      1 dårörtens
      1 däröver
     20 därpå
      1 darra
      1 darrighet
      6 darrningar
     26 därtill
      1 därunder
      1 därute
      5 därutöver
     16 därvid
      3 därvidlag
      2 darwin
      1 darwinismen
      2 darwinistisk
      1 darwins
      2 dasami
      1 dash
      1 dashi
      1 dashibuljongen
      1 dashkosten
      1 dashmodellen
      1 dashstudien
      3 dåsighet
      2 dåsigheten
      3 dat
     39 data
      3 databas
      4 databasen
      1 datablad
      1 databussar
      2 datachips
      1 datahantering
      1 dataingångar
      1 datainsamlingstiden
      1 datainspektionen
      1 datalagringssystem
      1 datamängden
      1 datamängder
      1 datan
      1 datanätverk
      1 dataprogram
      1 dataskärmar
      1 datera
      1 daterad
      2 daterade
      1 daterades
      1 daterar
      1 dateras
      1 daterat
      2 daterats
      1 datering
      5 dåtida
      7 dåtidens
     14 dator
      1 datoranvändning
      1 datorarbete
      1 datorbaserad
      2 datorbaserade
      1 datorbearbetas
      1 datorbildskärmar
      1 datorchip
      8 datorer
      1 datorerna
      1 datorernas
      1 datorgenererad
      2 datorkommunikation
      1 datorledning
      1 datorminne
      1 datormodeller
      1 datormus
      5 datorn
      2 datorövervakning
      4 datorprogram
      1 datorprogramvara
      4 datorskärm
      6 datorspel
      1 datorspelande
      1 datorspelen
      1 datorspelsfusk
      1 datorstödda
      4 datorsystem
      1 datorsystemet
      1 datortomograf
      3 datortomografen
     33 datortomografi
      1 datortomografibilder
      1 datortomografiguidad
      1 datortomografisk
      3 datortomografiundersökning
      1 datorutveckling
      8 datum
      3 datumet
      4 datummärkning
      1 datummärkningen
      2 datummärkta
      1 datura
      1 dauvers
      8 dåvarande
      1 davatarer
      1 davbildning
     10 david
      1 davidii
      1 davids
      3 davidson
      2 davis
      3 davy
      1 davyum
      1 day
     26 db
     10 dba
      2 dbild
      1 dbilder
      1 dbp
      1 dbrist
      1 dbt
      1 dbvärdena
      1 dc
      1 dcc
      2 dcd
      1 dckopplad
      1 dcläge
      2 dcs
      1 [dcs]
      2 dd
      1 ddd
      2 ddeprenyl
      7 ddimer
      1 ddimerkoncentrationen
      2 dds
     21 ddt
      1 ddts
      1 ddttoleranta
   5282 de
      2 dead
      1 deamidering
      1 deaminerar
      4 dean
      3 death
      1 deathrelated
      1 deaubonne
     15 debatt
     15 debatten
      1 debatter
      1 debatterad
      2 debatterades
      2 debatterar
      2 debatteras
      2 debatterat
      1 debatterats
      1 debranchingenzym
      1 debriefing
      9 debut
      1 debutålder
      1 debutåldern
      4 debuten
      6 debutera
      1 debuterade
      2 debuterande
     10 debuterar
      1 debuterat
      1 debutsymptomen
      1 debutsymtom
      2 debyescherrermetoden
      2 dec
      1 decade
      1 decades
      1 decalvans
     27 december
     18 decennier
     12 decennierna
      1 decenniernas
      3 decenniet
      5 decennium
      3 decentraliserad
      1 decentraliserat
      2 decety
      3 decibel
      1 decimalskala
      1 decimerades
      3 decimeter
      1 decimeterbred
      1 decimeters
      1 decinficering
      1 decipiens
      1 deckare
      1 decokten
      1 décolletage
      1 décolleter
      1 decompression
      1 decreased
      1 decumbens
      2 dederich
      1 dedicerat
      1 dee
      4 deep
      1 deer
      1 deet
      2 def
     20 defekt
      2 defekta
      9 defekten
     11 defekter
      1 defekterna
      1 defense
      2 deferens
      2 defiant
      1 defibrillator
      5 defibrillatorer
      2 defibrillera
      9 defibrillering
      1 defibrilleringsbar
      1 defibrilleringsbara
      4 deficit
      1 deficits
     11 definiera
      2 definierad
     11 definierade
      4 definierades
     18 definierar
     69 definieras
     13 definierat
      1 definierats
     61 definition
     19 definitionen
      2 definitionens
     20 definitioner
      3 definitionerna
      4 definitionsmässigt
      7 definitiv
      2 definitiva
      1 definitivsvar
      8 definitivt
      3 deformation
      1 deformationen
      2 deformerad
      2 deformerade
      1 deformerar
      3 deformeras
      1 deformeringen
      2 deformitet
      1 deformiteten
      1 deformiteter
      1 defosforyleringar
      4 deg
      2 degen
      7 degeneration
      3 degenerativa
      1 degenerera
      1 degenererade
      3 degenereras
      1 degenererats
      1 degeneres
      1 degig
      1 degranulera
      1 degranuleras
      1 degranulering
      2 degree
      1 dehumanisering
      1 dehydratiseras
      1 dehydratiseringsmedel
      1 dehydrerad
     11 dehydrering
      1 dehydroaripiprazol
      4 dehydroepiandrosteron
      1 dehydroepiandrosteronsulfat
      1 dehydrogenas
      1 dehydrogenation
      1 dehydrohalogeneras
      1 deimos
      1 déja
      2 dejoderas
      1 dekalin
      1 dekarboxylering
      1 deklaration
      1 deklarationen
      1 deklarationer
      2 deklarera
      1 deklarerades
      2 deklarerar
      1 deklarerat
      1 deklination
      1 dekolletage
      1 dekompression
      3 dekompressionen
      1 dekompressionsbehandling
      6 dekompressionssjuka
      2 dekor
      1 dekorationer
      2 dekorativ
      2 dekorativa
      1 dekorera
      1 dekorerad
      1 dekorerade
      2 dekoreras
    636 del
     36 dela
      7 delad
     19 delade
      7 delades
      1 delaktig
      1 delaktiga
      8 delaktighet
      1 delaktigheten
      2 delaktigt
    344 delar
     19 delarna
      1 delarnas
    109 delas
      1 delaspekten
      7 delat
      1 delats
      1 delaware
      1 delayed
      1 delblad
      1 delbladen
      1 delbrueckii
      1 delegation
      1 delegationer
      1 delegera
      1 delegerar
      2 delegeras
      3 delegering
      2 delegeringen
      1 delement
    150 delen
      1 delens
      1 deleterat
      1 deletion
      1 delfiner
      1 delförening
      1 delfrukter
      1 delfunktioner
      1 delgrupperna
      1 delhi
      2 delhudsbrännskada
      1 delidentiteter
      1 delight
      3 delikatess
     29 delirium
      1 delkärnan
      5 delkärnor
      1 delkomponent
      2 delkomponenter
     11 delmål
      6 delning
      3 delningen
      1 delningsfasen
      1 delningsskåra
      1 delningstakt
      1 delnorticus
      1 delokaliserade
      1 delphi
      1 delphinium
      1 delrapporter
      1 delrapporterna
      1 delresultat
    248 dels
      1 delskalor
      5 delstater
      3 delstaterna
      1 delstation
      1 delstatlig
      1 delsymtom
      2 delsystem
     14 delta
      5 deltagande
      3 deltagare
      1 deltagaren
      1 deltagarens
      7 deltagarna
      1 deltakvadranten
      1 deltametrin
     18 deltar
      2 deltavåg
      5 deltog
      1 deltyp
     88 delvis
    394 dem
     39 demens
      1 demensdiagnos
      1 demensen
      1 demenser
      1 demensfall
      1 demenslika
      1 demenspatienter
      4 demenssjukdom
     11 demenssjukdomar
      1 demenssjukdomarna
      2 demenssjukdomen
      2 demenssymtom
      2 demenstillstånd
      1 demenstypen
      1 demensutredningarna
      1 demensvård
      1 dementa
      5 dementia
      1 demeure
      1 demineralisationshastighet
      2 demivegetarianer
      1 democratic
      1 demodexkvalster
      1 demodikos
      2 demografi
      4 demografiska
      2 demografiskt
      5 demokratiska
      6 demoner
      1 demonerna
      1 demoniskt
      1 demonologi
      2 demonstrationer
      1 demonstrera
      1 demonstrerar
      1 demonstrerat
      1 demontera
      4 demoskop
      1 demyelinisering
      1 demyeliseringssyndrom
   6623 den
      2 denatonium
      7 denatoniumbensoat
      1 denatoniumsackarid
      1 denatoniumsalter
      1 denaturera
      1 denaturerar
      1 denatureras
      1 denaturerat
      1 denaturerats
      1 denaturering
      2 denatureringsmedel
      3 dendrit
      2 dendritcellen
     15 dendriten
      2 dendritens
     17 dendriter
     12 dendriterna
      4 dendriternas
      4 dendritiska
      1 dendritstammen
      1 dendritstrukturen
      1 dendritstukturen
      1 dendritsynapserna
      3 dendrittaggar
      2 dendrittaggarna
      1 dendrittätheten
      1 dendrodendritiska
     60 dengue
      1 dengueblödarfeber
      5 denguechocksyndrom
      1 dengueepidemier
     45 denguefeber
      2 denguefebern
      1 denguesymptomen
      1 dengueutbrottet
      7 denguevirus
      9 dengueviruset
      1 denham
      1 denheter
      1 denis
    892 denna
      2 dennas
     25 denne
     20 dennes
      1 denneval
      2 dennis
      1 denovo
      1 densa
     18 densamma
     21 densitet
      6 densiteten
      2 density
      6 dental
      1 dentallösning
      4 dentata
      1 dentatus
      1 dentinet
      1 dentosal
      1 deoderantmärke
      5 deodorant
      2 deodoranten
      9 deodoranter
      1 deodorantkristall
      1 deodorantsprejen
      2 deoxihemoglobin
      1 deoxy
      1 deoxygenerat
      1 deoxyhemoglobin
      1 depå
      1 depåfett
      2 departement
      2 departementet
      1 departementschefen
      4 department
      1 dependability
      1 dependant
     20 depersonalisation
      2 depersonalisationen
      1 depersonalisations
      1 depersonalisationsstörning
      6 depersonalisationssyndrom
      1 depersonalistisk
      2 depilering
      1 depolarisaion
      2 depolarisation
      1 depolarisationen
      1 depolariserade
      1 depolariseras
      6 depolarisering
      3 depolariseringen
      3 deponeras
      1 deponeringsform
      2 deponi
      1 deponiavgifterna
      1 depoteffekt
      1 depressio
    179 depression
     16 depressionen
      1 depressionens
     39 depressioner
      2 depressionerna
      1 depressionsbehandling
      1 depressionsformen
      1 depressionsfrekvens
      1 depressionspsykos
      2 depressionstillstånd
      2 depressiv
      9 depressiva
      1 depressivitet
      6 deprimerad
     11 deprimerade
      2 deprivation
     14 der
    247 deras
     18 derealisation
      1 derealisationssyndrom
     12 derivat
      1 derivative
      1 dermahud
      1 dermalt
      1 dermatillofagi
     12 dermatillomani
      6 dermatit
      1 dermatitidis
      2 dermatitis
      1 dermatitiska
      2 dermatol
      3 dermatologer
      4 dermatologi
      1 dermatologia
      3 dermatom
      2 dermatomen
      3 dermatomyosit
      1 dermatophagoides
      1 dermatoskop
      1 dermatovenereologi
      1 dermed
      3 dermis
      1 dermoida
      1 dermoidcysta
      1 dermologie
      8 des
      6 desamma
      1 desaturation
      3 descartes
      1 descendens
      1 descenderat
      2 desensibilisera
      6 desensibilisering
      1 desensitization
      2 desfluran
      8 design
      2 designade
      2 designades
      1 designats
      2 designen
      1 designerdrog
      1 designers
      1 designföretag
      1 designkläder
     35 desinfektion
      2 desinfektionslösningar
     18 desinfektionsmedel
      2 desinfektionssprit
      3 desinficera
      2 desinficerande
      4 desinficeras
      1 desinficering
      1 desinficeringsmedel
      1 desintegrativ
      2 deskvamation
      1 deskvamativ
      1 desmeknoppsväxter
      1 desmetoxicurcumin
      2 desorganisation
      7 desorganiserat
     10 desorientering
      1 desorption
    461 dess
   1252 dessa
      6 dessas
      1 dessert
      1 dessertviner
      1 dessförinnan
    216 dessutom
      7 dessvärre
      4 destillation
      1 destillerar
      3 destilleras
      1 destillering
      1 destilleringen
      1 destination
      1 destinationen
      1 destinationens
      1 destinationsuppfödda
     53 desto
      1 destruera
      2 destrueras
      4 destruktion
      1 destruktionen
      1 destruktionsapparat
      1 destruktionsdrift
      3 destruktiv
      2 destruktiva
      1 destruktivitet
      1 destruktivt
   7959 det
      1 �det
      4 detalj
      1 detaljbearbetning
      1 detaljen
      7 detaljer
      3 detaljerad
      4 detaljerade
      1 detaljhandel
      1 detaljhandlare
      2 detaljkunskaper
      1 detaljnivå
      1 detaljseende
      1 detaljseendedetaljstyrning
      1 detaljstudier
      7 detektera
      1 detekterade
      3 detekterar
      3 detekteras
      1 detekterat
      2 detektering
      3 detektion
      2 detektor
      1 detektorer
      6 detektorn
      1 deten
      1 detergent
      3 detergenter
      1 determinism
     11 detet
      1 detonerar
      1 detoxeffekt
      1 detritus
     19 detsamma
   1787 detta
      1 dettadessa
      1 dettas
      1 dettaurvalökar
      1 dettweiler
      1 deus
      2 deusta
      1 deuteragonist
      1 deuteragonisten
      1 deutschen
      1 deux
      1 devalvering
      6 devanagari
      1 developed
      1 developmental
      7 dexametason
      1 dexamethasone
      6 dexamfetamin
      1 dexamfetaminsulfat
      1 dexedrine
      1 dexofen
      1 dexter
      6 dextran
      1 dextranmolekyl
      1 dextriner
      3 dextroamfetamin
      2 dextrometorfan
      3 dextropropoxifen
      2 dextros
      1 dfilm
      4 dglukos
      1 �dglukos
      7 dhatu
     11 dhea
      1 dhenin
      3 dhfr
      6 dht
      2 dhumapana
      1 dhumpana
      2 dhupa
      1 dhyana
      2 di
      1 dia
      1 diabaínein
    166 diabetes
      1 diabetesen
      1 diabetesform
      3 diabeteskoma
      2 diabetesnefropati
      1 diabetespatienter
      2 diabetessjuka
      1 diabetessjuksköterskor
     19 diabetiker
      1 diachrolux
      1 diadem
      3 diafragma
      4 diafragmabråck
      3 diafragmamuskeln
      3 diafragman
      1 diafragmans
      2 diagfragmabråck
    274 diagnos
      1 diagnosbegrepp
      1 diagnosbeskrivningar
    150 diagnosen
      1 diagnosenabscesser
      1 diagnosens
     55 diagnoser
      1 diagnoseras
      1 diagnosering
     15 diagnoserna
      1 diagnosformer
      1 diagnosgrupper
      1 diagnosindelning
      1 diagnosinstrument
      1 diagnosis
      1 diagnosiska
      1 diagnosklassificering
      1 diagnoskod
      1 diagnoskoder
      1 diagnoskravet
      6 diagnoskriterier
      5 diagnoskriterierna
      4 diagnosmanual
      4 diagnosmanualen
      6 diagnosmanualer
      2 diagnosmanualerna
      1 diagnosmässigt
      1 diagnosmetod
      1 diagnosmetoden
      1 diagnosmetoder
      1 diagnossättet
      1 diagnosställning
      2 diagnossystem
      1 diagnosteknik
     10 diagnostic
      7 diagnosticera
      3 diagnosticerade
      2 diagnosticerar
     22 diagnosticeras
      1 diagnosticerats
      6 diagnosticering
      2 diagnosticeringen
      1 diagnosticeringskriterier
      1 diagnosticers
      1 diagnostiesera
     60 diagnostik
      8 diagnostiken
      4 diagnostillfället
     48 diagnostisera
      4 diagnostiserad
     11 diagnostiserade
      2 diagnostiserades
      9 diagnostiserar
     31 diagnostiseras
      1 diagnostiserat
      6 diagnostiserats
      1 diagnostiserbart
     18 diagnostisering
      2 diagnostiseringen
      1 diagnostiseringsmanualen
     10 diagnostisk
     35 diagnostiska
      6 diagnostiskt
      1 diagonalen
      1 diagonser
      5 diagram
      1 diagrammet
      4 diakon
      1 diakonal
      2 dialektala
      1 dialektalt
      1 dialektform
      1 dialektisk
      4 dialog
      2 dialogen
      1 dialoger
      1 dialogfilosofi
     13 dialys
      1 dialysapparater
      1 dialysator
      2 dialysatormembranet
      1 dialysatorn
      1 dialysavdelningen
      3 dialysbehandling
      1 dialysbehandlingen
      2 dialysen
      2 dialysera
      3 dialyserar
      1 dialyseras
      1 dialysfasen
      1 dialyskateter
      1 dialyskliniker
      1 dialyskoncentrat
      1 dialyskoncentratet
      1 dialyskrävande
      1 dialysmaskin
      1 dialysmaskinen
      1 dialysmembran
      1 dialysolyckan
      1 dialyspatienter
      1 dialysprocessen
      1 dialystillfälle
      2 dialysvätska
      4 dialysvätskan
      1 diamantförsedd
      1 diamantskallerorm
     42 diameter
      3 diametern
      1 diametrar
      1 diaminer
      1 diaminobensen
      1 diaminoxidas
      2 diamond
      1 dianoia
      2 diaphragman
     82 diarré
      1 diarreer
     17 diarréer
      2 diarréformen
      4 diarrén
      1 diarrér
      1 diarrésjukdom
      2 diarrésjukdomar
      1 diárroia
      1 diarylketoner
      1 diaspor
      2 diasporer
      1 diasporor
      1 diatermi
      3 diaton
      1 diaz
      2 diazepam
      1 dibutylftalat
      1 dibutyltenn
      2 dic
      1 dicentra
      2 dichelobacter
      1 dicke
      1 dickens
      1 dickinson
      3 dicom
      1 dictionnaire
      1 dicumarol
      3 did
      5 die
      1 dielstanus
      2 diemba
      1 diencephalon
     27 diet
      1 dietary
      1 dietbehandling
      1 dietbehandlingen
     28 dieten
      1 dietens
      6 dieter
      4 dieterna
      1 dieternas
      1 dietetic
      1 dietetik
      1 dietetiken
      1 diethylstilbestrol
      1 dietics
      1 dietik
      1 dietiskt
      8 dietist
      2 dietisten
      4 dietister
      1 dietitians
      1 dietplanen
      1 dietplaner
      1 dietrich
      8 dietylenglykol
      1 dietylenglykolen
      2 dietyleter
      1 dietylkarbamazin
      2 dietylstilbestrol
      1 dieu
      1 difenyl
      1 difenylketon
      1 differemtiis
      1 differences
      1 differentiade
      1 differential
      5 differentialdiagnos
      1 differentialdiagnosen
      8 differentialdiagnoser
      1 differentialdiagnostik
      1 differentialdiagnostiken
      1 differentialdiagnostiska
      1 differentialdiagostiska
      4 differentiating
      1 differentiell
      1 differentiera
      3 differentierad
      3 differentierade
      2 differentierar
      1 differentieras
      5 differentiering
      1 diffraktionsgitter
      1 diffraktionsmönster
      1 diffraktionsmönstret
      2 diffraktionspunkterna
      1 diffundera
      7 diffunderar
      9 diffus
     15 diffusa
     18 diffusion
      1 diffusiontack
      1 diffust
      2 diflucan
      1 difluordiklormetan
      6 difluorklormetan
      1 difluorklormetann
      7 difteri
      1 difteritoxinet
      1 difteroida
      9 dig
      1 digenea
      1 digeorge
      1 digeorges
     23 digerdöden
      4 digerdödens
      1 digestion
      1 digestionsenzym
      1 digestionsenzymet
      1 digestionskanalen
      1 digestionssystemet
      1 digher
      6 digital
     20 digitala
      1 digitale
      1 digitalform
      1 digitalin
      6 digitalis
      1 digitaliserar
      1 digitalisliknande
      1 digitalissläktet
      6 digitalt
      1 digitatus
      1 digiti
      1 digitoxin
      1 digitus
      1 dignostisering
      1 dihalometanen
      1 dihydroergocristine
      1 dihydroergocryptinmesilat
      1 dihydroergokorninmesylat
      1 dihydroergotamin
      1 dihydrofolat
      1 dihydrofolatreduktas
      3 dihydropteroatsyntetas
      4 dihydrotestosteron
      1 �dihydrotestosteron
      1 dihydroxibensen
      1 dihydroxifenoler
      1 dihydroxybensen
      1 dijodtyrosin
      1 dike
      2 diken
      1 dikeskanter
      2 diklofenak
      1 diklofenakpreparat
      1 dikloracetater
      1 dikloracetatjonen
      4 diklorättiksyra
      1 diklordifenyltrikloretan
      1 diklorkarben
      2 diklormetan
      1 diklorpropan
      2 dikotomi
      1 dikotomin
      4 dikt
      1 diktaturer
      1 dikten
      1 dikter
      1 dikteras
      1 dikterats
      1 diktform
      2 diktning
      1 diktsamlingen
      2 dikumarol
      2 dikväveoxid
      2 dilatera
      1 dilaterade
      1 dilaterar
      1 dilatering
      1 dilavore
      1 dilemma
      2 dille
      1 dilthey
      1 dimensioer
      3 dimension
      1 dimensionell
      1 dimensionen
     11 dimensioner
      1 dimensionerat
      1 dimensionerna
      1 dimensionslösa
      1 dimer
      2 dimeren
      1 dimeriseras
      1 dimerisering
      2 dimetylsulfat
      1 dimetylxantin
      1 dimidiatum
      1 diminutiv
      2 dimma
      1 dimmig
      2 dimsyn
      7 din
      1 dinga
      1 dingla
      1 dinitrofenol
      1 dioder
      1 diodorus
      3 dioica
      1 diol
      1 dionysiska
      1 dionysius
      1 dionysos
      2 dioptric
      2 dioptrier
      1 dioptriskt
      1 dior
      1 diorit
      2 diors
      2 dioskorides
      1 dioxidiamidoarsenobensol
      2 dioxin
      6 dioxiner
      1 dioxoantracen
      1 diphtheriae
      1 diploblastiska
      5 diploid
      7 diploida
      2 diplokocker
      1 diplom
      1 diplomatin
      1 diplomerad
      3 diplomerade
      1 dipsia
      2 dipsomani
      1 dipsomania
      1 dipsos
      1 diptera
      1 diptericin
      1 diras
      1 dire
      1 direction
      1 directthe
    215 direkt
     22 direkta
      1 direktion
     11 direktiv
      4 direktivet
      1 direktivets
     11 direktkontakt
      2 direktör
      2 direktörerna
      1 direktöversättning
      3 direktsända
      3 direktstimulerande
      1 direkttransfusion
      1 direktuppkopplade
      2 direktverkande
      1 diresorcin
      1 dirigerar
      3 disc
     10 disciplin
      2 disciplinen
      8 discipliner
      1 disciplinnämnd
      1 disco
      2 discovery
     20 disease
      6 diseases
      1 diseaseviruset
      5 disk
      4 diska
      1 diskanthörselnedsättning
      1 diskantljud
      5 diskar
      1 diskarna
      4 diskas
      1 diskbalja
      2 diskbaljor
      3 diskbänk
      1 diskbänkar
      1 diskbänken
      1 diskborste
      3 diskbråck
      4 disken
      7 diskgodset
      1 diskhandduk
      4 diskho
      2 diskit
      1 diskläge
      9 diskmaskin
     10 diskmaskinen
      1 diskmaskinens
      3 diskmaskiner
      1 diskmaskinerna
      1 diskmaskins
      7 diskmedel
      1 diskmedlet
      7 diskning
      3 diskningen
      1 diskogena
      1 diskonteras
      2 diskontering
      1 diskontinuerlig
      1 diskontinuerliga
      1 diskordanta
      1 diskotek
      1 diskoteksbesök
      1 diskrepans
      2 diskret
      1 diskreta
      1 diskriminerande
      1 diskrimineras
      5 diskriminering
      1 diskrimineringen
      1 diskställ
      1 disksvampar
      1 disktiden
      1 disktrasa
      2 disktrasor
      1 diskurser
      1 diskurserna
      2 diskus
     10 diskussion
      3 diskussionen
      3 diskussioner
      1 diskussionerna
      9 diskutera
      3 diskuterades
      4 diskuterar
      9 diskuteras
      3 diskuterat
      4 diskuterats
      1 diskuterbart
      1 diskvatten
      1 dislokaliseras
     14 disorder
     13 disorders
      1 dispalur
      2 dispens
      1 dispensärdistrikt
      1 dispensärer
      2 dispenserna
      2 dispergerade
      1 dispergeringsmedel
      3 display
      1 displayen
      2 dispositionsrätt
      1 disproportionalitet
      1 disputerade
      1 disputerat
      1 dispyter
      1 disse
      1 dissekerande
      3 dissektion
      3 dissektioner
      2 disseminerad
      1 dissertation
      1 dissident
      1 dissidenter
      3 dissociation
      1 dissociationen
      1 dissociationskurva
      1 dissociationsteori
      1 dissociationstillstånd
     14 dissociativ
     14 dissociativa
      1 dissociativt
      4 dissocierar
      1 distala
      3 distalt
      1 distance
      7 distans
      1 distanserar
      1 distansering
      1 distansutbildning
      1 distemper
      1 distinct
      3 distinkt
      2 distinkta
      5 distinktion
      1 distinktionen
      1 distortion
      2 distrahera
      1 distraherande
      2 distraheras
      1 distrahering
      1 distraktionsfri
      4 distress
      3 distresser
      1 distribuera
      4 distribueras
      2 distribution
      2 distributionen
      1 distributionskedjan
      1 distributionsledningar
      1 distributionsnät
      1 distributionsnätverk
      3 distributionssystem
      1 distributionsvolymen
      1 distributiv
      1 distributörer
      1 distributors
      2 distrikt
      1 distriktet
      1 distriktsbarnmorskor
      2 distriktsläkare
      2 distriktsnivå
      2 distriktssköterskor
     31 dit
      1 dithörande
      1 ditionit
      1 ditomyldijodid
      8 ditt
      5 dittills
      1 diuresi
      2 diuretika
      1 divalenta
      1 divergensen
      1 divergerande
     24 diverse
      2 diversilobum
      1 diversitet
      1 divertiklar
      1 divertikulos
      1 dividerad
      1 dividerades
      2 divideras
      3 dividerat
      1 dividing
      1 divigel
      1 divinorum
      1 division
      2 divisioner
      1 divisum
      1 divoire
      1 dizziness
      1 djävlar
      3 djävulen
      1 djävulens
      1 djävulsris
      1 djävulssopp
      1 djingis
     41 djup
     28 djupa
      1 djupalexi
      1 djupandning
     38 djupare
      1 djupaste
      1 djupavspänning
      3 djupberusning
      1 djupberusningens
      3 djupet
      1 djupfryst
      1 djupfrysta
      1 djupgående
      1 djuphavet
      1 djuphavsarter
      1 djupinvasiv
      1 djupliggande
      1 djupmätare
      1 djuppsykologi
      1 djupröda
      3 djupseende
      1 djupsömnen
      1 djupsömnsterapi
     25 djupt
    306 djur
      2 djurart
     18 djurarter
      1 djuraveln
      2 djurben
      1 djurbesättningar
      1 djurbestånd
      1 djurbon
      3 djurceller
     24 djuren
      9 djurens
      2 djurepitel
     40 djuret
      4 djurets
      1 djurexperiment
      1 djurfobiker
      2 djurfoder
     38 djurförsök
      1 djurförsöksetisk
      2 djurförsöksetiska
      2 djurförsöksstatistik
      1 djurfri
      1 djurgruppen
      1 djurhållare
      2 djurhållning
      2 djurhälsa
      1 djurhälsopersonal
      2 djurhannar
      1 djurindustri
      1 djurindustrin
      4 djurkadaver
      1 djurkliniker
      1 djurkontroller
      1 djurkroppar
      1 djurkroppen
      2 djurliv
      3 djurlöss
      5 djurlössen
      1 djurmodell
      4 djurpark
      2 djurparken
      5 djurparker
      1 djurparksbesökare
      1 djurplågeri
      2 djurpopulation
      1 djurrättsaktivister
      1 djurrättsorganisationen
      4 djurriket
      7 djurs
      1 djursjukdom
      1 djursjukhus
      1 djursjukskötare
      1 djursjukskötarprogrammet
      1 djursjukvård
      3 djursjukvårdare
      1 djursjukvårdaren
      1 djursjukvårdarlinjen
      1 djursjukvårdarnas
      1 djursjukvårdarprogrammet
      2 djursjukvården
      2 djurskötare
      1 djurskötaren
      2 djurskydd
      1 djurskyddet
      1 djurskyddslagstiftning
      1 djurskyddsmyndigheten
      1 djurskyddsorganisationer
      1 djurskyltar
      1 djurslag
      2 djurstudier
      1 djurtandvård
      1 djurtarmar
      4 djurtester
      1 djurtesterna
      1 djurvård
      2 djurvårdare
      1 djurvården
      2 djurvärlden
      2 dkf
      1 dkraftplattor
      1 dkupa
      2 dl
      3 dlaktat
      1 dlaktatet
      1 dlaktatrest
      1 dlb
      1 dl�tokoferol
      1 dm
      1 dmard
      1 dmitrij
      1 dmodellen
      1 dmsa
      1 dmscds
      2 dmt
      2 dn
     39 dna
      1 dnaanalys
      1 dnabaserade
      1 dnabildningen
      1 dnachips
      2 dnaforskning
      2 dnagyras
      2 dnamolekylen
      1 dnamolekyler
      1 dnamolekylerna
      1 dnanivå
      1 dnareplikation
      1 dnasekvenser
      2 dnasträngar
      1 dnasyntesen
      2 dnat
      1 dnateknik
      1 dnatest
      1 dnavaccin
      1 dnavirus
      1 dnp
      1 do
     34 dö
      1 dobson
      2 docent
      1 docetaxel
    938 dock
      2 docka
      1 dockhem
      1 dockögon
      1 dockorna
      1 dockteater
      3 doctor
     78 död
     94 döda
      2 dödad
      8 dödade
      7 dödades
      4 dödande
     29 dödar
      1 dödare
      8 dödas
      7 dödat
      3 dödats
      1 dödboksnotiser
     80 döden
      1 dödens
      1 dödenupplevelser
      6 dödfödda
      1 dödföds
      2 dödfödsel
      1 dödförklaring
      3 dödfött
     55 dödlig
     19 dödliga
      2 dödligaste
     36 dödlighet
     38 dödligheten
      1 dödlighetsprocenten
      1 dödlighetssiffrorna
     12 dödligt
      1 döds
      1 dödsÅngset
      1 dödsbegreppet
      2 dödsbo
      1 dödsbringande
      2 dödsdömde
      1 dödsdriften
    110 dödsfall
      1 dödsfallår
      8 dödsfallen
      7 dödsfallet
      1 dödsfallssiffran
      1 dödsguden
      3 dödshjälp
      1 dödskalle
      1 dödskriterier
      2 dödsoffer
      1 dödsoffren
      1 dödsögonblicket
      2 dödsolyckor
      1 dödsolyckorna
      9 dödsorsak
     12 dödsorsaken
      4 dödsorsaker
      9 dödsorsakerna
      1 dödspulver
      4 dödsriket
      1 dödsrisken
      1 dödssiffrorna
     10 dödsstraff
      3 dödsstraffet
      3 dödstal
      2 dödstalen
      1 dödstalet
      1 dody
      3 döende
     20 doft
      1 dofta
      1 doftämne
      2 doftämnen
      3 doftande
      3 doftar
      4 doften
      2 dofter
      1 doftflaggan
      1 doftlös
      1 doftlösa
     58 dog
      2 dogonfolket
      1 dogs
      1 doidge
      1 doing
      6 dök
      8 doktor
      1 doktorerade
      1 doktorn
      1 doktorsavhandling
      1 doktorsavhandlingen
      3 doktorsexamen
      1 doktorstitel
      1 doktrin
      4 dokument
      3 dokumentär
      1 dokumentärfilmen
     12 dokumentation
      1 dokumentationen
      1 dokumentationsarbete
      3 dokumentera
      5 dokumenterad
     22 dokumenterade
      3 dokumenterar
      9 dokumenteras
     11 dokumenterat
      9 dokumenterats
      1 dokumentering
      1 dokumenteringen
      2 dokumentförstörare
      4 dold
      2 dolda
      1 dolere
      1 dolikocefal
     10 dölja
      1 döljas
      4 döljer
      3 döljs
      1 dolk
      1 doll
     17 dollar
      2 dolomit
      1 dolomite
      1 dolor
      1 dolorosa
      4 dom
      1 döma
      2 domagk
      2 dömande
      1 domänen
      1 domäner
      1 domar
      1 domarboken
      1 domare
      1 domaren
      1 domarna
      1 domarnas
      3 dömas
      1 dömda
      6 dömde
      8 dömdes
      2 domen
      1 domens
      1 domesticerade
      1 domesticerat
      1 domestikationen
      2 dominans
      1 dominansen
      1 dominanskolumner
      7 dominant
      2 dominanta
      2 dominera
      3 dominerade
      1 dominerades
     19 dominerande
     14 dominerar
      7 domineras
      3 dominerat
      1 dominerats
      1 dominianus
      1 domkyrkan
      1 domnade
      3 domning
      8 domningar
      1 domningssymptomen
      1 döms
      1 domslut
      5 domstol
      2 domstolar
      1 domstolarna
      2 domstolen
      1 domstolens
      1 domstolsprövning
      3 dömts
      1 don
      2 donald
      2 donationer
      8 donator
      1 donatorbakterien
      6 donatorer
      1 donatorn
      1 donatorns
      1 donatorsperma
      3 donepezil
      2 donera
      2 donerad
      2 donerade
      3 donerar
      3 doneras
      1 donezepil
      1 donna
      1 donné
      2 dop
      1 dopamet
     19 dopamin
      1 dopaminagonist
      2 dopaminagonister
      2 dopaminaktiviteten
      1 dopaminåterupptag
      1 dopaminbetahydroxylas
      1 dopaminer
      3 dopaminerg
      4 dopaminerga
      1 dopaminet
      2 dopaminets
      1 dopaminförande
      1 dopaminfrisättande
      2 dopaminhypotesen
      1 dopaminkatabolitiska
      1 dopaminnivåerna
      2 dopaminreceptorer
      3 dopaminreceptorerna
      1 dopaminsignaleringen
      1 dopaminstabiliserare
      1 dopamintransportören
      1 dopaminutsöndringen
      1 döparen
      1 dopas
      1 dopbäcken
      6 doping
      1 dopingklassat
      2 dopingpreparat
      4 dopning
      2 dopningsklassat
      1 dopningspreparat
      1 dopningsskandaler
      2 dopp
      1 doppa
      3 doppade
      1 doppades
      2 doppas
      3 doppler
      2 dopplerteknik
      1 doppskor
      3 döpte
      1 doptique
      1 döpts
     85 dör
      1 dorn
      1 dörr
      5 dörrar
      1 dörren
      1 dörrhandtag
      2 dörrklocka
      1 dörrvakt
      1 dörrvakter
      1 dörrvakts
      3 dorsalis
      1 dorsalklipp
      1 dorsalrot
      1 dorsalsnitt
      1 dortmund
     73 dos
      1 dosa
      1 dosapotek
      1 dosberoende
      4 dose
     22 dosen
      1 dosens
      1 dosepainting
     72 doser
      1 dosera
      1 doserade
      2 doserar
      7 dosering
      1 doseringarna
      5 doseringen
      1 doseringsfärdiga
      1 doseringsform
      1 doseringsslarv
      4 doserna
      1 doses
      1 dosfritt
      2 doshas
      1 dosimetri
      1 doskonformitet
      1 dosoberoende
      1 dosområde
      1 dospåsar
      1 dosplan
      2 dosplanen
      1 dosplaner
      1 dosplaneringspersonal
      1 dosplaneringsprogram
      1 dosplaneringsprogrammet
      4 dosplaneringssystem
      1 dosplaneringssystemet
      1 dosplanerna
      1 dospotenta
     14 dosrat
      1 dosreduktion
      2 dosrespons
      3 dosresponskurva
      1 dosresponskurvor
      1 dosresponssamband
     20 dött
      9 dotter
      6 dotterbolag
      1 dotterbolagen
      1 dotterbolaget
      4 dotterceller
      2 dottercellerna
      1 dottercellernas
      3 dottern
      1 dotterplantor
      1 dottersvulst
      2 dottersvulster
      4 dottertaxa
      4 döttrar
      4 double
      1 doubt
      1 douche
      2 douglas
      2 doula
      6 döv
     15 döva
      1 dövahörselskadade
      1 dovare
      1 dövas
      4 dövblind
     13 dövblinda
      1 dövblindas
      3 dövblindblivna
      1 dövblinde
      3 dövblindfödda
      8 dövblindhet
      1 dövblindheten
      1 dövblindtolkar
      1 dövblint
     11 dövhet
      2 dövstumma
      1 dövt
      1 dowicide
     10 downs
      1 doxorubicin
      1 doxycyclin
      9 doxycyklin
      2 dpotenser
      1 dqdq
     30 dr
     56 dra
     51 drabba
     25 drabbad
    279 drabbade
     40 drabbades
    155 drabbar
    281 drabbas
      9 drabbat
     74 drabbats
      3 drack
      2 dracunculus
     41 drag
      1 dragbo
      2 dragen
      1 dräger
      1 dragera
      1 drages
      2 dragit
      1 dragkamp
      1 dragkedja
      1 drägligt
      4 dragning
      2 dragningskraft
      1 dragok
      1 dragon
      1 dragsjuka
      1 drakar
      2 drake
      1 drakhuvuden
      1 drakhuvudet
      1 dräkt
      2 dräkten
      3 dräkter
      3 dräktiga
      1 dräktighet
      4 dräktigheten
      1 dräktjackor
      2 drama
      1 dramafilmen
      1 dramaserie
      1 dramaserien
      2 dramat
     10 dramatisk
      5 dramatiska
      8 dramatiskt
      1 drän
      3 dränage
      1 dränaget
      4 dränera
      1 dränerar
      7 dräneras
      1 dränering
      1 dräneringen
      1 dräneringsanordning
      1 dräneringskateter
      1 dräng
      2 dränka
      1 dränkning
      1 dränseras
      3 dråp
      1 dråpare
      1 dräpt
     44 drar
     45 dras
      1 drastica
      1 drastisk
      5 drastiska
      9 drastiskt
      1 dravyaguna
      1 dream
      1 dreaming
      1 dreceptorer
      1 dresden
      1 dressad
      1 dressing
      7 drev
      4 drevs
      2 dri
     42 dricka
      3 drickande
      1 drickas
      1 drickbart
     13 dricker
      1 drickes
      4 dricks
      1 dricksglas
     17 dricksvatten
      1 dricksvattenproduktion
      6 dricksvattnet
      5 drift
      4 driften
     10 drifter
      3 drifterna
      2 driftparametrar
      2 driftsäkerhet
      1 driftsäkerhetsmåttet
      1 driftskostnaderna
      1 driftsliv
      1 driftteori
      1 drig
      1 drill
      1 drink
      1 drinkar
      1 drinkarna
      2 drinking
      1 drinkingwater
     11 driva
      1 drivas
      4 driven
     17 driver
      4 drivit
      2 drivits
      2 drivkraft
      1 drivkraften
      1 drivkrafter
      1 drivkrafterna
      2 drivmedel
      1 drivremmar
      1 drivrutiner
     14 drivs
      2 drivsystemet
      1 drivtryck
      1 drnovšek
     35 drog
      1 droganvändarna
      9 droganvändning
      1 drogarbete
      2 drogavvänjning
      3 drogberoende
      3 drogbruk
      1 drogbrukaren
      2 drogbrukarna
     24 drogen
      2 drogens
     94 droger
      4 drogerna
      1 drogförebyggande
      3 drogförgiftning
      2 drogframkallade
      2 drogfrihet
      2 drogintag
      1 drogkonsumenten
      6 drogkonsumenter
      2 drogkonsumtion
      1 drogkonventioner
      9 drogmissbruk
      1 drogmissbrukare
      1 drogpåverkade
      1 drogpåverkan
      1 drogpåverkat
      4 drogpolitik
      3 drogpolitiken
      1 drogrelaterade
      2 drogrus
     13 drogs
      1 drogsmugglaren
      3 drogtest
      2 drogtester
      1 drogtrafiken
     15 drogutlöst
      9 drogutlösta
      1 dröj
      5 dröja
      3 dröjde
      2 dröjer
      1 dröjsmål
      6 dröm
      1 drömfarare
      1 drömforskning
      1 drömframkallande
      1 dröminnehåll
      1 drömlika
      1 drömliknande
      1 drömmande
     19 drömmar
      1 drömmare
      1 drömmaren
      3 drömmarna
      5 drömmen
      6 drömmer
      1 drömsekvensen
      5 drömsömn
      1 drömsömnen
      1 drömsömnstadiet
      1 drömteori
      1 drömterapi
      2 drömtydning
      2 drömvärlden
      1 drönare
      1 drop
      6 dropp
      5 droppa
      1 droppades
      1 droppande
     17 droppar
      1 droppas
      2 droppe
      2 droppen
      1 droppform
      3 droppfot
      4 droppsmitta
      1 dror
      9 drottning
      1 drottningar
      1 drottningen
      1 drottningsubstans
      1 drs
      1 drsp
      4 druckit
      1 druckits
      9 drug
      1 drugbank
      6 drugs
      2 drunkenness
      1 drunkna
      1 drunknade
     11 drunkning
      1 drunkningskänslor
      1 drunkningsolyckor
      1 druvan
      1 druvans
      5 druvbörd
      2 druvfläder
      1 druvhinna
      2 druvhinnan
      4 druvhinneinflammation
      1 druvklasar
      1 druvklase
      1 druvliknande
      1 druvmusten
      2 druvor
      2 druvorna
      5 druvsocker
      3 druvsorter
      1 drycj
     20 dryck
      5 drycken
     17 drycker
      1 dryckers
      1 dryckeskärl
      1 dryfta
      3 dryg
      4 dryga
     43 drygt
      2 ds
      4 dserin
     17 dsm
      3 dsmiii
      2 dsmiiir
     30 dsmiv
      7 dsmivtr
      1 dsmmanualen
      1 dsms
      1 dsmsystemet
      4 dsmv
      1 dsmvtr
      2 dsps
      1 dsrna
      1 dss
      3 dst
      1 dstruktur
      1 dstrukturen
     10 dt
      1 dtenterografi
      1 dtpa
     60 du
      1 duac
      1 dualismen
      1 dualister
      1 dualistisk
      1 dubach
      2 dubbdäck
      8 dubbel
      4 dubbelbefruktning
      2 dubbelbindning
      3 dubbelbindningar
      2 dubbelbindningen
      1 dubbelblind
      2 dubbelblinda
      1 dubbelblindplacebokontrollerad
      2 dubbeldiagnos
      1 dubbeldiagnosen
      1 dubbeldiagnoser
      2 dubbellager
      1 dubbelmask
      1 dubbelriktad
      1 dubbelsaltet
      4 dubbelsidig
      1 dubbelsidigt
      2 dubbelskikt
      1 dubbelskiktet
      1 dubbelslag
      2 dubbelslipade
      1 dubbelsträngat
     14 dubbelt
      1 dubbeltecknas
      1 dubbelverkande
     11 dubbla
      1 dubblerade
      1 dubblerat
      1 dubius
      1 dubrovnik
      1 duchennes
      1 duct
     16 ductus
      1 dudaim
      1 dudley
      1 duell
      1 duffyblodgruppssystemet
      1 duglighet
      2 duk
      1 duka
      3 dukar
      1 dukarna
      2 duke
      2 dukemetoden
      1 dukes
      1 dukoral
      4 duktala
      1 duktig
      1 duktilitet
      1 duktus
      1 dulcamar�
      4 dulcamara
      1 dulcis
      2 dumas
      1 dumbe
      1 dumheter
      1 dumpade
      1 dumpades
      1 duncan
      2 duncans
      1 dunckers
      1 dunhårig
      1 dunhåriga
      2 dunkel
      4 dunkerque
      1 dunkningar
      1 dunkuddar
      1 dunn
      1 dunsta
      1 dunstar
      6 duodeni
      1 duodenojejunalis
     13 duodenum
      1 duplex
      1 duplexteknik
      1 dupliceras
      4 dupont
      1 durasäcken
      1 durat
      1 dürers
      1 during
      1 durissus
      2 durkheim
      1 durklopp
      1 durra
      1 durrakäppar
     14 dusch
      2 duscha
      1 duschaggregat
      1 duschandes
      6 duschar
      1 duschdraperi
      1 duschen
      1 duschgolv
      1 duschkabin
      1 duschkabinen
      2 duschning
      3 dussin
      1 dussintal
      1 duvbröst
      1 dux
      2 dvala
      2 dvärg
      4 dvärgar
      3 dvärgbandmask
      1 dvärgbandmasken
      1 dvärgelefanten
      1 dvärgkastning
      1 dvärgtyper
     12 dvärgväxt
      1 dvdn
      1 dverklighet
      1 dviruset
      8 dvitamin
      2 dvitaminbrist
      1 dvitaminer
      1 dvitaminmetabolismen
    117 dvs
      6 dvt
      1 dw
      1 dy
      1 dygderna
     67 dygn
      2 dygnen
     27 dygnet
      1 dygnetruntlinser
      1 dygnetruntrådgivning
      1 dygnsproduktion
      9 dygnsrytm
      4 dygnsrytmen
      1 dygnsrytmsjukdom
      1 dygnsurinmängd
      8 dyk
     15 dyka
      2 dykapparat
      1 dykapparaten
      1 dykardatordykarklockor
      1 dykardräkt
      1 dykardräkten
      1 dykardräkterna
     10 dykare
      7 dykaren
      1 dykares
      1 dykarklocka
      1 dykarklockor
      1 dykarklockorna
      1 dykarkomplikationer
      1 dykarloppor
      3 dykarna
     11 dykarsjuka
      2 dykarsjukan
      1 dykarskador
      1 dykartermer
      1 dykdator
      9 dyker
      1 dykmedicin
     11 dykning
      1 dykningar
      1 dykningens
      1 dykningfara
      1 dykningsolyckor
      1 dykorganisationer
      2 dykreflexen
      1 dykt
      1 dyktabeller
      3 dylik
      4 dylika
     14 dylikt
      1 dyna
      1 dynamic
      1 dynamik
      2 dynamiken
      1 dynamisering
      7 dynamisk
      5 dynamiska
      1 dynamo
      1 dynamometamorfos
      1 dynan
      1 dynod
      2 dynoden
      2 dynoder
      2 dynodkedjan
      1 dynvial
      5 dyr
      6 dyra
     13 dyrare
      2 dyraste
      1 dyrbar
      2 dyrbara
      1 dyrbaraste
      1 dyrkad
      1 dyrkade
      2 dyrkan
      8 dyrt
      6 dys
      1 dysa
      8 dysartri
      1 dysartrin
      5 dysbarism
      1 dyscalculia
      6 dysenteri
      1 dysenteriae
      1 dysenteribakterier
     25 dysfagi
      1 dysfagin
      3 dysfasi
      4 dysfoni
      2 dysfori
      3 dysforisk
      1 dysfunction
     50 dysfunktion
      3 dysfunktionell
      2 dysfunktionella
      1 dysfunktionellt
      2 dysfunktioner
      1 dysgalactiae
      1 dysgeusi
      2 dysgrafi
      1 dysgrafin
      1 dysgrammatism
      1 dysgraphia
     10 dyskalkyli
      3 dyskinesi
      1 dyskinesierna
      1 dyslektikerns
      1 dyslektiska
      1 dyslektiske
     22 dyslexi
      1 dyslexia
      1 dyslexidiagnos
      1 dyslexiförbundet
      1 dyslexiföreningen
      9 dysmeli
      1 dysmeliskadorna
      2 dysmenorré
      1 dysmnesi
     12 dysmorfofobi
      1 dysmorfofobisk
      1 dysmorphic
      8 dyspareuni
      1 dysphoros
      9 dysplasi
      2 dysplasia
      3 dysplasier
      1 dysplasierna
      1 dysplastisk
      7 dyspné
      1 dysport
      1 dyspraktisk
      2 dyspraxi
      1 dysprosodi
      1 dyssomni
      1 dyster
      1 dysterhet
      2 dyston
      2 dystoni
      1 dystonier
      1 dystra
      1 dystrofin
      3 dystymi
      1 dystymier
      4 dysuri
      1 dyvelsträck
     99 e
      1 ea
      2 eagt
      1 eagtackrediterat
      1 eanox
      2 eap
      3 ear
      1 earle
      2 early
      1 east
      2 eastman
      1 eat
      3 eata
      1 eatas
      3 eau
      1 ebbe
      1 ebenezer
      1 ebenholts
      1 eberhard
      6 ebers
      1 eberspapyrusen
      1 eboga
     30 ebola
      9 ebolafeber
      1 ebolafebern
      1 ebolafloden
      1 ebolainfekterad
      1 ebolainfektioner
      1 ebolautbrott
      1 ebolautbrotten
      2 ebolautbrottet
      1 ebolavironets
     16 ebolavirus
      9 ebolaviruset
      2 ebolavirusets
      2 ebonit
     19 ebrt
      1 ebrtbehandlingen
      1 ebulus
      1 ebv
      1 ec
      1 ecc
      1 eccegodkänt
      1 ecdc
      1 echa
      2 echelon
      1 echinaceas
      1 echinaceatillskott
      5 echinococcos
      2 echinococcus
      4 echinokockinfektion
      1 echis
      1 echo
      1 echolalia
      1 eciwobaserad
      1 eck
      1 eckinokockos
      1 ecnn
      1 École
      6 ecoli
      1 ecology
      1 ecosoc
      2 ecstasy
      1 ecstasypiller
     21 ect
      7 ectbehandling
      3 ectbehandlingar
      2 ectropion
      1 ectserie
      4 ecuador
      1 ecuadorianska
      7 ed
      3 edema
      1 edematosa
      1 eder
      1 ederöversättning
      1 edet
      1 edguy
      1 edifact
      3 edinburgh
      3 edith
      3 edition
      1 edlén
      2 edler
      1 edmond
      1 edmund
      4 edoperioden
      1 Édouard
      1 edra
      1 edta
      1 eduard
      1 eduardo
      7 education
      1 educations
      1 edvard
      9 edward
      2 edwards
      1 edwardsson
      3 edwin
      1 edzard
      3 ee
     21 eeg
      1 eegmätning
      1 eegmätningar
      1 eegundersökningen
      1 eelementet
      1 efedrin
      2 effect
      1 effectivness
      1 effects
      1 effekivt
    302 effekt
     88 effekten
    116 effekter
     49 effekterna
     67 effektiv
     57 effektiva
     17 effektivare
      4 effektivast
      3 effektivaste
      1 effektiviseras
     16 effektivitet
      6 effektiviteten
     94 effektivt
      1 effektivtatt
      1 effektorcell
      1 effektpedal
      2 effektstyrka
      1 effektstyrkan
      2 efferenta
      1 efflux
      1 effluxfunktion
      1 effluxprotein
      1 effusion
   1453 efter
     25 efteråt
      1 efterbearbetning
      2 efterbehandlas
      1 efterbehandling
      3 efterbliven
      1 efterblödning
     10 efterföljande
      6 efterföljare
      1 efterföljarstater
      2 efterföljd
      4 efterföljs
      1 efterföljt
      4 efterförloppet
      1 efterforskningar
     12 efterfrågan
      3 efterfrågas
     21 efterhand
      1 efterhärmar
      1 efterkoncentrationen
      1 efterkontroll
      1 efterkrigsbarnen
      2 efterladdaren
      4 efterladdning
      2 efterladdningssystem
      1 efterladdningsteknik
      1 efterladdningsutrustning
      1 efterlämnade
      1 efterleden
      1 efterledet
      1 efterlevande
      1 efterlevandes
      1 efterlevas
      1 efterlevnad
      3 efterlevs
      3 efterlikna
      1 efterliknade
      1 efterliv
      1 efterloppet
      1 efterlysningen
      2 eftermiddagen
      1 efternamn
      1 eftersedimentering
      1 eftersläpning
      1 eftersmak
      1 eftersök
      1 eftersökta
    742 eftersom
      2 eftersträvade
      4 eftersträvas
      1 eftersträvat
      1 eftersvettning
      1 eftertänksamhet
      1 efterträdde
      1 efterträddes
      1 efterträder
      2 eftertraktade
      1 eftertraktades
      1 eftertraktat
      1 eftervakuum
      1 eftervårdsprogram
      1 eftervärlden
      1 efterverkningarna
     12 eg
      2 egas
      3 egdomstolen
    118 egen
      1 egenart
      2 egenartad
      1 egenarten
      3 egenbehandling
      1 egenbilden
      1 egenbrus
     10 egendom
      1 egendomliga
      1 egenföretagare
      1 egenförsörjning
      1 egenhändigt
      1 egenhet
      1 egenheter
      2 egenkontroll
      1 egenmakt
      1 egennamn
      1 egenrehabilitering
     22 egenskap
     13 egenskapen
    149 egenskaper
     16 egenskaperna
      1 egentillverkat
     14 egentlig
     18 egentliga
     53 egentligen
      3 egentligt
      7 egenvård
      2 egenvården
      1 egenvårdprimärvård
      1 egenvårdsbranschen
      1 egenvårdshäften
      1 egenvårdsråd
     45 eget
      1 egfr
      1 egfrinhibitorer
      1 eggar
    100 egna
      4 ego
      1 egodystona
      1 egodystoniska
      1 egoistiska
      1 egosyntona
      5 egot
     15 egypten
      2 egyptens
      1 egyptier
      5 egyptierna
      1 egyptiernakälla
      1 egyptiernas
      4 egyptisk
      9 egyptiska
      2 ehälsa
      1 ehinger
      2 ehlersdanlos
      1 ehrenkreuz
     11 ehrlich
      1 ehrlichhata
      7 ehrlichios
      2 ehrlichs
      1 ei
      1 eikosanoider
      1 eiloés
      2 einar
      3 eindhoven
      1 eine
      1 einecs
      1 einer
      1 einsiedeln
      1 einstein
      2 einthoven
      2 einthovens
      1 eisacktal
      1 eisenberg
      1 eisenbergs
      1 eitrem
    143 ej
      3 ejakulatet
     13 ejakulation
      7 ejakulationen
      1 ejakulationens
      1 ejakulatorisk
      1 ejakulatoriska
      1 ejakulerade
      1 ejakulerar
      1 ejektionsfraktion
      1 ek
      1 eka
      1 ekdysteron
      1 ekerliknande
     20 ekg
      1 ekganalyser
      1 ekgapparat
      1 ekgapparaten
      1 ekgapparatens
      1 ekgapparater
      2 ekgförändringar
      1 ekgförändringarna
      1 ekgkurva
      2 ekgmätning
      2 ekgt
      1 ekgtester
      1 ekgundersökning
      1 ekgundersökningar
      1 ekgutseendet
      4 eklampsi
      2 eklampsiutveckling
      1 eklöf
      2 eklund
      1 eko
      2 ekofeminism
      1 ekofeminismen
      2 ekokardiografen
      9 ekokardiografi
      2 ekokardiografins
      1 ekokardiografiutrustningar
      1 ekokardiogram
      1 ekokardiogrammet
      4 ekolali
      1 ekoliknande
      1 ekolod
      9 ekologi
      2 ekologin
      3 ekologisk
      2 ekologiska
      2 ekologiskt
      1 ekon
      1 ekonomerna
      9 ekonomi
      1 ekonomier
      3 ekonomin
      1 ekonomipriset
     11 ekonomisk
     39 ekonomiska
     11 ekonomiskt
      1 ekorrar
      1 ekorre
      1 ekosymtom
      6 ekosystem
     15 ekr
     34 eksem
      1 eksematös
      5 eksemet
      1 eksemlika
      1 eksemliknande
      1 eksempatienter
      1 ekström
      1 ektallskogar
      2 ektoderm
      3 ektome
      2 ektoparasit
      3 ektoparasiter
      3 ektopisk
      1 ektopiska
      1 ektoterm
      1 ekvation
      3 ekvationen
      1 ekvatorialregionen
      3 ekvatorn
      1 ekvilibrium
      5 ekvivalent
      4 ekvivalenta
      6 el
      1 elaffärer
     21 elakartad
     18 elakartade
      2 elakartat
      2 elakt
      1 elakupunktur
      2 elallergi
      1 elapider
      1 elapiders
      6 elasticitet
      2 elasticiteten
      2 elastin
      5 elastisk
      9 elastiska
      7 elastiskt
      2 elastografi
      1 elavskärmande
      1 elbehandling
      2 elbehandlingar
      1 elbow
      1 elbs
      1 elbsreaktionen
      1 elcentraler
      4 elchocker
      1 elchockpistoler
     20 eld
      1 eldades
      2 eldar
      1 eldas
      1 elddon
      4 elden
      1 eldfasta
      1 eldhärden
      2 eldmakande
      1 eldning
      1 eldningsmaterial
      1 eldriven
      2 eldrivna
      1 eldslåga
      2 eldslagning
      2 eldsoffer
      1 eldstad
      1 eldstaden
      1 eldstunga
      1 eldsvåda
      1 eldsvådor
      2 eldticka
      4 eldtickan
      1 eldtorn
      1 eleanor
      2 electric
      2 electrical
      2 electroconvulsive
      1 electronic
      6 electronics
      1 electrospray
      1 electuarium
      3 elefant
      2 elefanten
      4 elefanter
      7 elefantiasis
      1 elefantlusen
      1 elefantmannen
      1 elefantnäbbmusen
      1 elegans
      1 elegant
      3 eleganta
      1 elektomagnetisk
      7 elektricitet
      2 elektriker
     41 elektrisk
     79 elektriska
     20 elektriskt
      7 elektrod
      4 elektroden
     20 elektroder
     10 elektroderna
      2 elektrodernas
      1 elektrodplacering
      1 elektrodplaceringen
      1 elektrodrad
      1 elektrodstimulering
      2 elektroencefalografi
      1 elektroencefalogram
      1 elektrofil
      3 elektrofilter
      1 elektroforetiska
      1 elektrofysiologi
      1 elektrofysiologisk
      1 elektrokardiografi
      1 elektrokardiogram
      3 elektrokemisk
      1 elektrokemiska
      3 elektrokonvulsiv
      4 elektrolys
      1 elektrolysen
      3 elektrolyt
      1 elektrolytbalans
      5 elektrolytbalansen
      4 elektrolyten
     15 elektrolyter
      1 elektrolyterna
      1 elektrolytisk
      1 elektrolytiska
      1 elektrolytkoncentrationerna
      2 elektrolytlösningar
      1 elektrolytnivåer
      1 elektrolytproduktion
      1 elektrolytrubbningen
     13 elektromagnetisk
     16 elektromagnetiska
      1 elektromekanisk
      1 elektrometer
      1 elektromyograf
      1 elektromyografen
      3 elektromyografi
      1 elektromyogram
      4 elektron
      1 elektrondensitetskarta
      1 elektrondensitetskartan
      2 elektronens
     12 elektroner
      4 elektronerna
      4 elektroneurografi
      5 elektronik
      1 elektronikfackhandeln
      1 elektronikindustrin
      1 elektronikkonstruktioner
      1 elektronikprylar
      1 elektroniktillverkare
      1 elektroniktillverkarna
      8 elektronisk
      9 elektroniska
      2 elektroniskt
      1 elektronmikrograf
      4 elektronmikroskop
      1 elektronmikroskopet
      1 elektronrör
      1 elektronsprejjonisering
      1 elektronstråle
      4 elektronstrålen
      1 elektronstrålning
      1 elektrontransporten
      4 elektrontransportkedjan
      1 elektrontransportproteiner
      1 elektrookulografi
      2 elektrostatisk
      3 elektrostatiska
      1 elektrotekniken
     11 element
      1 elementär
      1 elementära
      1 elementärt
      7 elementen
      1 elenergi
      2 eleonora
      1 elephantis
      5 elev
      1 elevated
      2 elevens
     16 elever
      1 elevernas
      2 elfenben
      1 elfte
      1 elgard
      2 elgitarr
      1 eliade
      1 elimination
      1 eliminationsförsök
      2 eliminationshalveringstid
      1 eliminationskost
      1 eliminationsreaktion
     16 eliminera
      1 eliminerades
      3 eliminerar
      5 elimineras
      1 eliminerat
      2 eliminerats
      3 eliminering
      1 elin
      6 elinder
      1 eliot
      7 elisa
      1 elisabetanska
      1 elisabeth
      1 elisany
      1 elisatest
      4 elit
      3 eliten
      2 elitidrottare
      1 elitträning
      1 elittrupper
      5 elizabeth
      1 elkabel
      1 elkablar
      1 elkänslighet
      1 elkoagulation
      1 elkostnad
      1 elkraft
      1 elledning
      2 ellen
   5895 eller
      1 ellermaskar
      1 ellerrimantadin
      3 ellipse
      8 elliptiska
      1 elliptiskt
      1 elmotordrivet
      1 elmotorer
      1 elmotorerna
      1 elongatus
      1 elöverkänslig
      6 elöverkänsliga
      3 elöverkänsligas
     15 elöverkänslighet
      1 elproduktion
      1 elradiatorer
      7 elsanering
      2 elsevier
      1 elstandard
      1 elstatus
      1 elstötar
      4 eltandborstar
      5 eltandborste
      1 eltandborsten
      1 eltandborstens
      1 elton
      1 eluttag
     10 elva
      1 elvahundratalet
      3 elvanse
      1 elver
      2 em
      2 ema
      1 email
      6 emalj
      5 emaljen
      1 emaljens
      1 emaljerad
      1 emaljöga
      1 emaljytan
      1 emanerar
      1 emanuel
      1 emanuella
      7 emboli
      1 emboliserar
      2 embolisk
      1 emboliska
      1 embolism
      2 embolus
      8 embryo
      1 embryoblaster
      1 embryodonation
      1 embryofyter
      1 embryogenes
      2 embryogenesen
      1 embryologiska
      2 embryon
      2 embryonal
      3 embryonala
      1 embryonalt
      2 embryoperioden
     15 embryot
      1 embryotfostretbarnet
      4 embryots
      1 emc
      6 emdr
      3 emedan
      1 emedicine
      5 emellan
      5 emellanåt
    106 emellertid
      1 emergency
      1 emerson
      1 emetica
      2 emetika
      2 emfnet
      2 emfysem
     20 emg
      1 emi
      2 emigranter
      1 Émile
      1 emilie
      1 emilio
      2 emiscanner
      4 emission
      1 emissioner
      1 emissions
      1 emissionsspektrum
      1 emit
      1 emitteras
      1 emlakräm
      2 emma
      1 emo
      1 emorroides
     61 emot
      7 emotionell
     14 emotionella
     11 emotionellt
      3 emotioner
      1 emotions
      1 emotionspsykologi
      1 empasote
      3 empaten
      1 empater
      1 empatheia
      1 empathic
      3 empathy
     55 empati
      1 empatibegreppet
      1 empatibegreppets
      1 empatiforskning
      1 empatiforskningen
      1 empatilös
      1 empatilöshet
      6 empatisk
      6 empatiska
      1 empatiskt
      1 empatisystem
      3 empatisystemet
      1 empatiträning
      3 empiri
      4 empirisk
      2 empiriska
      5 empiriskt
      1 emplastrum
      1 employment
      7 empyem
      1 ems
      1 emsömn
      2 emulgera
      1 emulgerar
      1 emulsin
      6 emulsion
      1 emulsionen
      4 emulsioner
      1 emycin
  13767 en
    100 ena
      4 enades
      1 enäggssyskon
      1 enäggstolvlingar
      1 enäggstvåtuslingar
      2 enäggstvilling
      7 enäggstvillingar
      1 enäggstvillingen
      1 enahanda
      1 enan
      1 enantiomerer
      3 enantiomererna
      1 enarmade
      1 enas
      2 enastående
      1 enbär
    142 enbart
      1 enbaspolymorfier
      1 enbrel
      9 encefalit
      1 encefaliter
      2 encefalitvirus
      4 encefalopati
     10 encelliga
      1 encelligt
      2 encephalitis
      1 enco
      2 encyklopedin
    129 enda
      1 endags
      1 endagslinser
      1 endangered
    441 endast
      3 endemi
      3 endemicum
      1 endemios
     11 endemisk
      4 endemiska
      2 endemiskt
      8 endera
      1 endexpiratory
      1 endimensionella
      1 endimensionellt
      1 endo
      1 endocyterar
      6 endocytos
      1 endoderm
      1 endodermal
      1 endodonti
      1 endodontin
      1 endodontisk
      2 endofenotyp
      1 endofenotyper
      4 endogen
      4 endogena
      1 endogent
      1 endokardiet
     11 endokardit
      2 endokardium
      1 endokardos
     12 endokrin
     68 endokrina
      1 endokrinkirurgi
      1 endokrinologen
      2 endokrinologer
      7 endokrinologi
      1 endokrinologin
      1 endokrinologisk
      7 endokrint
      4 endometriet
      1 endometriomas
     21 endometrios
      1 endometrioscystor
      1 endometriosdrabbade
      3 endometriosen
      1 endometriospatienter
      1 endometriosveckan
      1 endometrit
      3 endoplasmatiska
      1 endorfin
      4 endorfiner
      1 endorsement
      1 endoscopy
      4 endoskop
      3 endoskopet
      5 endoskopi
      3 endoskopisk
      1 endoskopiska
      1 endosomerna
      2 endosomet
      1 endospermet
      1 endostatin
      1 endostin
      2 endosulfan
      7 endotel
     20 endotelceller
      9 endotelcellerna
      2 endotelcellernas
      1 endotelet
      1 endotelin
      3 endotelium
      1 endotelprogenitorceller
      1 endoterm
      1 endothelial
      1 endotoxin
      9 endotoxiner
      1 endotoxinerna
      1 endotoxinhaltiga
      1 endotoxisk
      2 endotrachealtub
      2 endotrakealtub
      1 endotrakealtuben
      1 endotrakealtuber
      1 endovaskulärt
      1 endrokrin
      6 eneg
      2 enegmätningar
      1 enegmätningarna
      1 enegundersökning
      1 energeidrycker
      1 energetik
     72 energi
      1 energiapparater
      1 energiatomära
      1 energibegrepp
      2 energibegreppet
      5 energibehov
      1 energibehovet
      1 energibesparande
      1 energibrist
      2 energicentra
      1 energidrycken
      1 energidrycker
      1 energieffektiv
      8 energier
      1 energifält
      1 energiförbränningen
      5 energiförbrukning
      1 energiförbrukningen
      1 energiförlust
      1 energiförråd
      1 energiförsörjningsmekanismer
      1 energifunktion
      1 energiindustrin
      1 energiinnehåll
      4 energiinnehållet
      5 energiintag
      4 energikälla
      2 energikällor
      1 energikick
      6 energikrävande
      1 energilager
      1 energilöshet
      2 energimängd
      1 energimängden
      2 energimärkning
      4 energimärkningen
      1 energimässiga
      1 energimässigt
      1 energimedicinska
      1 energimetabolismen
      1 energimyndigheten
      8 energin
      1 energinivåer
      1 energiöverskottet
      1 energiprincipen
      1 energiproduktion
      2 energireserv
      1 energireserver
      2 energirika
      3 energisk
      1 energiska
      1 energiskt
      1 energismart
      2 energisnåla
      1 energisnålt
      1 energisystem
      1 energitäthet
      1 energitillförsel
      1 energityperna
      1 energiunderskott
      1 energiutbytet
      1 energiutvinningen
      1 energivärde
      1 energivärdet
      1 enfluran
      1 enforcement
      2 enformiga
      1 enformigt
      1 enfülhung
     17 eng
      7 engagemang
      1 engagement
      3 engagera
      1 engagerad
      3 engagerade
      1 engagerar
      5 engångs
      2 engångsbindor
      1 engångsblad
      2 engångsdos
      1 engångsdosering
      1 engångsföreteelse
      1 engångshanddukar
      1 engångshandskar
      1 engångskanyler
      1 engångskatetrar
      1 engångskonsumtion
      1 engångslinser
      1 engångsmaterial
      1 engångsmensskydd
      1 engångsmodell
      1 engångsprodukt
      1 engångsprodukter
      1 engångsskalpeller
      1 engångsskydd
      1 engångstratt
      2 engångsvarianter
      1 enge
     11 engelsk
    128 engelska
      9 engelskan
     12 engelskans
      8 engelske
      1 engelskspråkig
      3 engelskspråkiga
      4 engelskt
      1 engelsktalande
      1 engelsmän
      2 engelsmannen
      1 engelsmännen
      1 engelsmännens
      2 engineering
      2 engineers
     48 england
      1 englands
      1 englandslistan
      1 englewood
      1 english
      4 engström
      1 enhag
      1 enhancement
      9 enhet
     17 enheten
      6 enheter
      2 enheterml
      1 enheterna
      7 enhetlig
      4 enhetliga
      3 enhetligt
      1 enhetscell
      1 enhetscellen
      1 enhetsfel
      1 enhetsstruktur
      2 enhjärtbladiga
      1 enhörningshorn
      3 eniga
      1 enighet
      1 enigmatit
      1 enkät
      1 enkäten
      2 enkäter
      2 enkätstudie
      1 enkätundersökning
      2 enkefaliner
      1 enkefalinerga
     36 enkel
      1 enkelblommiga
      1 enkelinlärd
      1 enkelkedjigt
      2 enkelomättat
      2 enkelriktad
      3 enkelsidig
      1 enkelsträngad
      1 enkelsträngade
      3 enkelsträngat
     73 enkelt
     51 enkla
     44 enklare
      3 enklast
     14 enklaste
      2 enkoimesis
      6 enkönade
      2 enl
     19 enlighet
      1 enlighten
    482 enligt
      1 ennukleotider
      1 enol
      1 enorganismsmotståndskraft
     10 enorm
      8 enorma
      2 enormt
      1 enquireinquire
      1 enriched
      1 enrollerat
      1 enrummig
     45 ens
     10 ensam
      1 ensamarbete
      4 ensamhet
      1 ensamheten
     15 ensamma
      1 ensamme
      1 ensamrätt
      1 ensamrätten
      9 ensamstående
      8 ensamt
      1 ensessionsbehandling
      1 ensessionsbehandlingar
      1 ensessionsbehandlingen
     10 ensidig
      2 ensidiga
      3 ensidigt
      1 ensilage
      1 ensileringsmedel
      2 enskiktat
     18 enskild
     44 enskilda
     15 enskilde
      1 enskildes
     16 enskilt
      1 ensläktet
     49 enstaka
      1 enstyrke
      1 ental
      1 enteogen
      1 enteogener
      1 enteral
      1 enterica
      5 enteriska
      2 enteroartrit
      2 enterobacter
      3 enterobacteriaceae
      1 enterobius
      3 enterococcus
      2 enterocyter
      1 enterokocken
      7 enterokocker
      2 enterotoxin
      4 enterovirus
      1 enteroviruspcr
      1 enterprise
      1 entesalgier
      1 entesopatierna
      1 entoloma
      1 entolomataceae
      1 entonox
      2 entoptiska
      1 entre
      1 entré
      1 entréhallar
      2 entrén
      1 entreprenadavtal
      1 entreprenören
      1 entreprenörer
      1 entrévärd
      1 entropion
      1 entusiaster
      3 entydig
      2 entydiga
      2 entydigt
      1 enukleation
      9 enummer
      2 enumret
      1 enures
      1 enureslarm
      2 env
      1 envåningsbastun
      1 envar
      1 envärd
      3 envärda
      2 envärt
      1 envelope
      1 environ
      1 environmental
      1 envis
      1 envishet
      1 enwikipedia
     51 enzym
      8 enzymatiska
      1 enzymatiskt
      1 enzymbehandlingar
      1 enzymbrist
      2 enzymdefekter
      2 enzyme
      1 enzymelinked
      5 enzymen
     54 enzymer
      7 enzymerna
      1 enzymes
     57 enzymet
      1 enzymets
      1 enzymgift
      1 enzymkemi
      1 enzymkopplad
      2 enzymsystem
      1 enzymsystemet
      1 enzymteoretisk
      3 eog
      2 eoh
      1 eosin
      2 eosinofil
      3 eosinofiler
      1 ep
      3 epa
      1 epas
      1 epaxal
      1 ependymalceller
      1 epicondylit
      1 epicondylus
      1 epidauros
      1 epidaurus
     20 epidemi
      1 epidemic
      2 epidemica
      1 epidemicyklerna
     23 epidemier
      4 epidemierna
      1 epidemiliknande
     12 epidemin
      1 epidemiolgiska
      1 epidemiologer
     31 epidemiologi
      2 epidemiologin
      1 epidemiologins
      4 epidemiologisk
      5 epidemiologiska
      1 epidemisjukhus
      4 epidemisk
      7 epidemiska
      1 epidemivåg
      2 epidermal
      1 epidermiphyton
      2 epidermis
      1 epidermophyton
      2 epididymis
      3 epididymit
      1 epiduo
      4 epiduralbedövning
      1 epifora
      4 epifysen
      1 epifysens
      2 epiglottis
      1 epigyn
      1 epikardiet
      2 epikardium
      1 epiklorhydrin
      1 epikondyl
      2 epikondylit
      1 epilambanein
      2 epilator
      1 epilatorer
      1 epilatorn
     53 epilepsi
      1 epilepsia
      4 epilepsianfall
      1 epilepsianfallens
      1 epilepsiframkallande
      1 epilepsikirurgi
      1 epilepsikirurgiskt
      2 epilepsiliknande
      1 epilepsimedicin
      1 epilepsimediciner
      4 epilepsin
      1 epilepsisjukdom
      1 epilepticus
      4 epileptiker
      2 epileptisk
     24 epileptiska
      7 epileptiskt
      2 epilering
      1 epinefrin
      1 epipharynx
      2 episk
      2 episod
      1 episoden
     11 episoder
      1 episoderna
      1 episodisk
      4 episodiska
      1 epispadi
      1 epistaxis
      1 episteme
      7 epitel
      1 epitelbeklädnaden
      1 epitelcell
     15 epitelceller
      5 epitelcellerna
      1 epitelcellernas
      4 epitelet
      1 epitelets
      1 epitellager
      1 epitelmuskelceller
      1 epiteloida
      1 epiteloidceller
      1 epitelyta
      1 epitet
      5 epithalamus
      1 epitlet
      4 epitoper
      1 epitoperna
      2 epizooti
      1 epizootilagen
      1 epizootilagstiftningen
      1 epizootiologi
      7 epo
      1 epodopning
      2 epok
      1 epoken
      1 epoker
      1 epomops
      1 Époque
      1 epost
      1 eposta
      1 epostmeddelanden
      2 epoxi
      1 epoxider
      1 epoxidgrupp
      1 epoxietan
      1 epoxiharts
      1 epoxilim
      1 epoxiplast
      1 epoxiplaster
      1 epsteinbarr
      3 epsteinbarrvirus
      1 ept
      3 eq
      1 equal
      2 equality
      1 equestre
      1 equi
      2 equina
      2 equinovarus
      1 equiperdum
      1 equivalent
      5 er
      1 eradictation
      2 eran
      3 eranthis
      3 erasmus
      1 erbach
      1 erbb
      7 erbjöd
      4 erbjöds
      6 erbjuda
      1 erbjudande
      2 erbjudanden
     12 erbjudas
     24 erbjuder
      2 erbjudit
      1 erbjudits
     21 erbjuds
      1 erc
      1 [erc]
      2 ercp
      1 ercs
      1 erdmann
      1 erecta
      2 erection
      1 eregerade
     37 erektil
      1 erektila
     33 erektion
     11 erektionen
      1 erektionens
      4 erektioner
      2 erektionerna
      3 erektionsförmågan
      1 erektionsperioder
      3 erektionsproblem
      1 erektionsproblemen
      1 erektionsstarten
      1 erektionsstörning
      1 erektionssvikt
      1 erektionssvikten
      1 eremitkräftor
      5 erfara
      1 erfaranhet
      4 erfaren
     25 erfarenhet
      5 erfarenheten
     27 erfarenheter
      1 erfarenheterna
      1 erfarenhetsmässig
      1 erfarit
      1 erfarna
      1 erforderliga
      2 erforderligt
      1 erfordliga
      1 erfordras
      1 ergenyl
      1 ergocornin
      1 ergocristin
      1 ergocryptin
      1 ergokalciferol
      1 ergoloidmesylat
      1 ergometrin
      1 ergometrintartrat
      2 ergon
     11 ergonomi
      1 ergonomisk
      1 ergonomiska
      1 ergonovin
      1 ergonovinmaleat
      3 ergotamin
      1 ergotamintartrat
      6 ergotism
      1 ergotoxinesilat
      1 ergotoxinfosfat
     14 erhålla
      1 erhållande
      5 erhållas
      1 erhållen
      5 erhåller
      4 erhålles
      3 erhållit
      4 erhållits
      1 erhållna
     12 erhålls
      1 erhart
      6 erhöll
      1 erhölls
      5 eric
      1 erich
      2 erickson
      1 ericksons
      1 ericsson
      1 ericssons
      3 erigerad
      1 erigeras
      2 erigerat
      1 erigeron
      5 erik
      1 erika
      3 erikson
      5 eriksson
      1 erikssons
      1 erinra
      1 erinus
      6 erkänd
      3 erkända
      5 erkände
      4 erkändes
      5 erkänna
      5 erkännande
      1 erkännanden
      3 erkännandet
      3 erkänner
      1 erkänns
      6 erkänt
      2 erland
      2 erlichia
      1 erlichiabakterien
      4 ernest
      3 ernst
      1 ernsthar
      1 eroderas
      1 erogena
      1 eros
      2 erosion
      1 erotica
      2 erotisk
      2 erotomani
      1 erövrare
      1 erövringen
      1 erowid
      1 erpositiv
      3 errector
      1 error
     10 ersatt
     25 ersätta
      1 ersättande
     13 ersättas
      7 ersatte
     14 ersätter
     12 ersattes
     18 ersättning
      1 ersättningar
      2 ersättningen
      1 ersättningmedel
      1 ersättningsföda
      1 ersättningsläkemedelsubstitution
      1 ersättningsmedel
      1 ersättningsrytm
      1 ersättningsrytmen
      1 ersättningsskyldig
     16 ersatts
     20 ersätts
      1 ersson
      1 ertharin
      3 ertms
      1 erudition
      2 erwin
      1 erwinia
      1 erygrocyterna
      1 eryhtrina
      1 erykah
      2 erysipelas
      1 erysiphales
      6 erytem
      2 erytema
      1 erytemen
      4 erythema
      3 erythematosus
      4 erytrocyt
      4 erytrocyten
      9 erytrocyter
      5 erytrocyterna
      1 erytrocyternas
      1 erytrocytkolinesterasaktivitet
      1 erytrocytkoncentrat
      1 erytrocytkoncentraten
      1 erytrocytproduktionen
      1 erytroida
      4 erytromycin
      2 erytropoes
      2 erytropoesen
      2 erytropoetin
      1 erytropoietinreceptorer
      1 erytros
      3 es
      1 esat
      6 esau
      1 esav
      1 esbittabletter
      4 esbl
      1 esblpositiva
      1 esblvarianter
      1 eschar
      9 escherichia
      1 eschscholtz
      1 eschscholzia
      1 esge
      2 esi
      1 esianvändas
      1 eskalerar
      1 eskulap
      2 esmark
      4 esofageal
      3 esofageala
      7 esofagus
      1 esofaguscancer
      3 esofagusvaricer
      1 esoterism
      3 espghan
      1 ess
      3 essay
      8 essel
      1 essels
      2 essenser
      3 essensoljor
      8 essentiell
      3 essentiella
      2 essentiellt
     13 essilor
      5 essilors
      1 esslingen
      1 establish
      2 esteban
      1 estelle
      3 ester
      1 esterbindningarna
      1 estermolekylerna
      1 estern
      1 esterreaktion
      1 estetikens
      7 estetisk
      7 estetiska
      4 estetiskt
      1 estimate
      1 estimating
      2 estimera
      3 estimeras
      1 estimerats
      3 estimering
      1 estland
      3 estradhypnos
      7 estrar
      1 esvl
      1 esyhaler
     35 et
      4 etablera
     10 etablerad
     27 etablerade
      8 etablerades
      2 etablerar
      2 etableras
      7 etablerat
      5 etablerats
      1 etablering
      2 etableringen
      1 etableringsrätten
      1 etablissemanget
      3 etac
      1 etambutol
      6 etan
      2 etanal
      6 etandiol
    102 etanol
      1 etanoldrift
      9 etanolen
      1 etanolförgiftning
      1 etanolmetaboliten
      1 etanolmolekylen
      1 etanolmolekyler
      1 etanolmotor
      2 etanols
      3 etansyra
      1 etansyran
      1 etappstoppen
     77 etc
      6 etcetera
      7 eten
      1 etenol
      1 etenoxid
     22 eter
      1 eteranestesi
      1 eterbedövning
      1 eterinhalationsnarkos
      1 eterisk
      9 eteriska
      1 eterkropp
      1 etern
     12 eternit
      1 eterniten
      1 eternitfabriken
      2 eternitplattan
      2 eternitplattor
      1 eternitskivor
      1 eternitskivorna
      1 etersövningen
      1 etest
      1 etex
      1 ethmoidale
      1 ethnocultural
      1 Étienne
      3 etik
      1 etiken
      1 etikens
      2 etikett
      2 etiketten
      2 etiketter
      1 etiketterad
      1 etiketterade
      1 etiketteras
      1 etinylöstradiol
     20 etiologi
      2 etiologier
      9 etiologin
      1 etiologisk
      1 etiologiskt
      4 etiopien
      1 etiopisk
      1 etiopiska
      4 etisk
      8 etiska
      8 etiskt
      3 etnicitet
      1 etniciteter
      2 etnisk
      9 etniska
      1 etnografen
      1 etnolog
      1 etnologin
      1 etnomedicin
      2 etologi
      1 etrar
      2 etsande
      2 etsning
   5643 ett
      1 [ett]
      1 ettan
      8 ettårig
      2 ettåriga
      1 ettårsåldern
      1 ettårsperspektivet
      1 ettårstudier
      1 ettbarnspolitik
      2 ettbetygskurserna
      1 ettbetygsnivån
      1 ettermyror
      1 etthundra
      1 etuiet
      3 etylacetat
      2 etylalkohol
      1 etylbensen
      1 etylbromid
      1 etylcellulosa
      1 etylcyanoakrylat
      1 etylcyanopropenoat
      1 etylen
      8 etylenglykol
      3 etylenglykolen
      1 etylenglykolförgiftning
      1 etylestern
      1 etyletanoat
      1 etylgrupp
      1 etylgrupper
      1 etylkatinon
      1 etylklorid
     30 etymologi
      2 etymologin
      1 etymologiskt
      1 etythrina
     41 eu
      1 euanpassad
      1 eublomman
      1 eucosmus
      2 eufemism
      1 eufemismen
      1 eufomani
      5 eufori
      2 euforin
      1 euforisk
      1 euforiska
      1 euforiskt
      1 euförordning
      4 eugen
      1 eugene
      1 eugenes
      7 eugenik
      4 eugeniken
      3 eugeniska
      1 eugenol
      1 eug�ne
      1 euhamn
      1 euinträdet
      1 eukalyptol
      6 eukaryota
      5 eukaryoter
      1 eukaryotiska
      5 eukommissionen
      1 eukommissionens
      1 eulagstiftning
      1 eulagstiftningens
      8 euländer
      1 euländers
      1 eumedborgare
      2 eumelanin
      1 eumoped
      2 eunivå
      2 eunucker
      2 euparlamentet
      1 eupatorium
      2 euphorbia
      2 euphorbiaceae
      1 eur
      3 eurasien
      1 eurekommendation
      5 euro
      3 eurobalis
      1 eurobalisen
      1 eurobaliser
      1 eurobaliserna
    197 europa
      1 europaea
      2 europafacket
      2 europakommissionens
      1 europakonventionen
      7 europaparlamentet
      3 europaparlamentets
      1 europarådet
      2 europarådets
     14 europas
      1 europastandard
      1 europe
     12 european
      1 europeanamerican
      1 européen
      8 européer
      3 européerna
      1 européernas
      1 européernordeuropéer
     11 europeisk
     78 europeiska
      2 europeiskt
      1 eurythmie
      9 eurytmi
      1 eurytmiensembler
     10 eurytmin
      4 eurytmins
      8 eus
      1 eustress
      1 eustressorer
      1 eutanasi
      1 euthyroid
      4 euthyroidsick
      1 eutrochium
      7 ev
      6 eva
      1 evacuare
      1 evakuerats
      2 evakuering
      2 evaluation
      1 evalueras
      1 evaluering
      1 evangelista
      1 evans
      1 evansi
      1 evaporering
      1 evar
      1 evd
      1 evenemang
      1 evenker
      1 evenki
     35 eventuell
     48 eventuella
     67 eventuellt
      1 evetuellt
      1 evf
      2 evidence
     11 evidens
      6 evidensbaserad
      1 evidensbaserade
      1 evidensbaserat
      1 evidensbasering
      4 evidensen
      2 evidensgrad
      1 evidensprövas
      1 evidensprövning
      1 evidensstudier
      1 evidensstyrka
      1 evidensundersökningen
      1 evig
      3 eviga
      1 evighet
      4 evigt
      1 evitamin
      1 evoked
      1 evoluon
      8 evolution
      7 evolutionär
      5 evolutionära
      8 evolutionärt
      1 evolutionella
      3 evolutionen
      1 evolutionistiska
      1 evolutionsbiologen
      1 evolutionsbiologi
      1 evolutionsforskning
      1 evolutionspsykologin
      1 evolutionsteori
      2 evolutionsteorin
      2 ewing
      9 ewings
      5 ewingsarkom
      1 ewloe
     99 ex
      1 exacerbation
     40 exakt
     23 exakta
      1 exalterad
     21 examen
      1 examensarbete
      1 examensnivå
      2 examensrätt
      1 examenstiteln
      1 examina
      1 examinan
      2 examination
      1 examinationer
      1 examinationsorganisationer
      2 examinerade
      2 examinerades
      1 examineradt
      1 examinerar
      1 examinerats
      1 exanthematicus
      1 exasperatum
      1 excavatum
      1 excellence
      1 excentricitet
      1 excentriker
      1 excentrisk
      1 excentriska
      1 excentriskhet
      1 excision
      1 excitatoriska
      2 excitera
      1 exciterad
      1 exciterar
      1 exciteras
      3 excitotoxicitet
      1 excitotoxologisk
      1 excrementerna
      5 executive
      2 exekutiv
      6 exekutiva
      1 exelon
      1 exemestan
   1331 exempel
    554 exempelvis
     27 exemplar
      2 exemplaren
      4 exemplaret
      3 exemplen
      1 exemplena
     11 exemplet
      2 exemplifierad
      1 exemplifierar
      4 exemplifieras
      1 exforge
      1 exhalterat
      1 exhibitionism
      8 existens
      7 existensen
      1 existensplanen
      3 existentiell
      4 existentiella
      4 existera
      5 existerade
     13 existerande
     37 existerar
      1 existerartroligtvis
      1 existerat
      1 existing
      1 exists
      1 exkluderade
      1 exkluderar
      1 exklusionskriterier
      2 exklusiv
      1 exklusivitet
      2 exklusivt
      1 exkret
      2 exkretion
      1 exocyterar
      8 exocytos
      1 exoftalmus
      1 exogena
      2 exogent
      5 exokrina
      6 exon
      1 exoner
      1 exorcism
      1 exoskelett
      2 exoterm
      1 exotiska
      1 exotiskt
      1 exotoxider
      3 exotoxin
      8 exotoxiner
      4 expandera
      1 expanderande
     12 expanderar
      2 expanderat
      1 expanderbara
      3 expansion
      1 expansionen
      1 expansionsplaner
      2 expedition
      1 expeditionen
      2 expeditioner
      1 expektoreras
      4 experience
     22 experiment
      5 experimentell
      3 experimentella
      5 experimentellt
      1 experimenten
      7 experimentera
      3 experimenterade
      1 experimentering
      3 experimentet
      1 experiments
      1 expert
      8 experter
      1 experterna
      1 expertgranskade
      1 expertgranskare
      1 expertgrupp
      1 expertgrupper
      1 experthjälp
      4 expertis
      1 expertsystemen
      1 expertutlåtanden
      1 expiratorisk
      4 expiratory
      1 explicita
      1 exploatera
      1 exploaterbart
      1 exploatering
      4 exploderar
      1 explorativ
      3 explorerande
      1 explosion
      3 explosionen
      1 explosionsartade
      2 explosionsartat
      2 explosiva
      3 explosivitet
      1 explosivt
      2 exponerad
      3 exponerade
      3 exponerades
      2 exponerar
     18 exponeras
      4 exponerats
     45 exponering
      3 exponeringar
     14 exponeringen
      1 exponeringsautomatik
      4 exponeringsbehandling
      1 exponeringskällan
      1 exponeringskategorierna
      1 exponeringsnivå
      1 exponeringsplatsen
      1 exponeringstabell
      1 exponeringstiden
      2 export
      2 exportera
      1 exporterade
      1 exportintäckter
      2 exportör
      1 exportunderskott
      1 exposed
      1 exposition
      1 exposure
      1 expressenjournalisten
      2 expression
      1 expressionsnivåer
      1 expressiva
      1 exspirationexhalation
      1 exsudativ
      3 extas
      1 extasiska
      1 extatisk
      1 extatiska
      1 extended
      1 extension
      1 extensioner
      1 extensivt
      1 extensorer
      9 extern
     36 externa
      1 externi
      3 externt
      1 externus
      1 extirpation
     82 extra
      2 extracellulär
      9 extracellulära
      1 extracellulärrummet
      4 extracellulärt
      1 extracellulärvätskan
      1 extracellullär
      1 extracellullära
      1 extracerebral
      1 extracerebralt
      1 extracorporeal
      1 extraction
      1 extractum
      5 extrafunktioner
      1 extrahepatiska
      3 extrahera
      2 extraherade
      2 extraheras
      1 extrakorporeal
      6 extrakt
      1 extrakten
      1 extraktet
      1 extraktion
      2 extraordinär
      1 extraordinära
      1 extrapontin
      5 extrapulmonell
      1 extrapunkter
      4 extrapyramidala
      3 extraslag
      1 extrautbildning
      1 extrauterin
      1 extrauterint
      1 extraventrikulärt
      1 extraversion
     25 extrem
     23 extrema
      1 extremely
      1 extremer
      1 extremfall
      3 extremitet
      3 extremiteten
     10 extremiteter
     14 extremiteterna
      3 extremitetsavledningar
      3 extremitetsavledningarna
      1 extremitetsförlusten
     53 extremt
      1 extremvärdet
      1 extrinsic
      1 extrinsikalt
      2 extrinsiska
      1 extroverta
      1 exudat
      5 eye
      1 eyelet
      1 eyeliner
      1 eyesyndromet
      1 eyre
      1 ezetrol
      1 ezhexadekadienol
     44 f
      2 �f
      1 fa
    665 få
      2 fabergé
      1 fabio
      1 fabrica
      1 fabricii
      8 fabrik
      3 fabrikat
      6 fabriken
      1 fabrikens
      4 fabriker
      1 fabriksframställda
      1 fabriksmässig
      1 fabriksmässigt
      1 fabrikstillverkade
      1 fäbroms
      3 face
      2 facebook
      1 facebookanvändare
      1 facebookvänner
      1 facettleder
      1 facettledsbesvär
      1 fachgebieten
      2 facialis
      1 facialisnerven
      3 facialispares
      1 facialisparese
      1 facialisparesen
      1 faciei
      1 facilities
      1 facing
      1 facitergium
      2 fack
      1 fackfolk
      2 fackförbund
      1 fackförening
      1 fackklubb
      1 fackkunskap
      2 fackla
      1 facklan
      1 fackliga
      1 fackligt
      1 fackmän
      1 fackområden
      1 fackorgan
      1 fackspråk
      1 facktidningar
      2 facs
      2 fact
      1 facto
     11 factor
      1 faculty
      9 fader
      4 fäder
     12 fadern
      1 fäderna
      1 faders
      1 fadersålder
      1 faderskap
      1 faderskapsundersökningar
      1 faecalis
      2 faeces
      1 faecesavgång
      2 faecium
      1 faengsel
      1 fåfänga
      8 fågel
      1 fågelägg
      3 fågelarter
      1 fågelbilharzia
      1 fågelbon
      1 fågelbröst
      1 fågeldjur
      6 fågelinfluensa
      3 fågelinfluensan
      1 fågellöss
      1 fågellössen
      2 fågeln
      1 fågelns
      1 fågelparasiter
      1 fågeluppfödare
     45 fåglar
      2 fåglarna
      1 fåglars
      2 fagocyter
      2 fagocytera
      1 fagocyterad
      1 fagocyterade
      2 fagocyterande
      2 fagocyteras
      1 fagocyterat
      3 fagocytos
      1 fagocytosen
      1 fagotten
      1 fagottens
      1 fåhr�us
      2 failure
      1 fair
      1 fairbairn
      1 fairly
      1 fak
      7 fakta
      1 faktaartiklar
      1 faktan
      1 fäktas
      3 faktisk
      9 faktiska
     35 faktiskt
      1 faktoid
     83 faktor
    179 faktorer
     13 faktorerna
      1 faktorernas
      1 faktorhalt
      2 faktorkoncentrat
     13 faktorn
     32 faktum
      1 faktureras
      3 fakultativt
      4 fakultet
      2 fakulteten
      1 fakulteterna
      1 falangen
      1 falciparum
    832 fall
     15 falla
      3 fälla
      1 fållade
      2 fällan
      1 fallande
      1 fallandesjuka
      1 fallandesot
      1 fällas
      1 fallbeskrivning
      2 fallbeskrivningar
      1 fällde
      2 fälldes
    111 fallen
      1 fallenhet
     46 faller
      2 fäller
     80 fallet
      1 fallets
      6 fallit
      1 fallkontrollstudie
      1 fall�kontrollstudie
      5 fällning
      1 fällningen
      1 fållor
      4 fällor
      1 fällorna
      1 fallosbärare
      1 fallossymbol
      2 fallossymboler
      2 fallrapporter
      1 fall�referentstudie
      1 fall�referentstudien
      7 fälls
      1 fällts
      6 falsett
      1 falsetten
      1 falsettsång
      2 falsettsångare
      1 falsifiera
      2 falsifierbar
      9 falsk
     15 falska
      8 falskt
      1 falso
     34 fält
      1 fälten
      7 fältet
      1 fältförhållanden
      1 fältförsök
      1 fältfritt
      1 fältherrarnas
      1 fältherren
      1 fälthygien
      1 fältläkare
      1 fältläkarreglementet
      1 fältmarskalken
      1 fältmössa
      1 fältmössor
      1 fälts
      1 fältsjukhus
      8 fältsjukvård
      6 fältskär
      1 fältskären
      1 fältskärer
      1 fältskärerna
      1 fältskog
      1 fältspatsgruva
      1 fältstyrkan
      1 fälttåg
      1 fältteori
      1 fältuniform
      1 falun
      1 falungongrörelsen
      1 famciklovir
     39 familj
      1 familjär
      4 familjebok
      1 familjefilmer
      1 familjehistoria
      1 familjehund
      1 familjeläkare
      2 familjeläkarmottagning
      3 familjelivet
      1 familjemässigt
      4 familjemedlem
      3 familjemedlemmar
      1 familjemedlemmarena
      1 familjemedlemmarna
      1 familjemedlems
    135 familjen
      3 familjens
      3 familjeplanering
      2 familjepolitik
     15 familjer
      1 familjerelationer
      1 familjerna
      1 familjernas
      1 familjestudier
      1 familjeterapi
      1 familjetragedi
      1 familjetvätteriet
      1 familjevänligt
      2 familjs
      2 fancy
      1 fåne
      3 fanerogamer
     11 fånga
      1 fångad
      1 fångade
     14 fångar
      1 fångaren
     11 fångas
      1 fångat
      1 fångats
     17 fängelse
      1 fängelseförbud
      2 fängelser
      2 fängelsestraff
      1 fängelsevåldtäkter
     17 fångenskap
      1 fangfolket
      1 fängslades
      1 fängslande
      1 fångsttrådar
      1 fångtransport
      1 fänkål
      1 fänkålsstänger
     44 fann
    131 fanns
      2 fänrikshjärtesläktet
      3 fantasi
      1 fantasieggande
      6 fantasier
      1 fantasiföreställningsförmåga
      1 fantasifulla
      1 fantasilösa
      1 fantasins
      1 fantastisk
      1 fantastiska
      1 fantastiskt
      1 fantasylitteraturen
      2 fantiserar
      2 fantomsmärta
     10 fao
      2 faos
      1 fap
      1 faq
     15 far
    784 får
     30 fara
      1 fårad
      1 faraday
     11 faran
      1 fåran
      1 farao
      1 faraonernas
      2 faraos
      1 fårbesättningen
      3 färd
      1 färdades
     14 färdas
      1 färdbroms
      1 färdhastighet
      5 färdig
     12 färdiga
      1 färdigberedd
      4 färdighet
      1 färdigheten
     12 färdigheter
      2 färdigheterna
      2 färdighetsträning
      1 färdigstädade
      1 färdigställandet
      1 färdigställer
      8 färdigt
      1 färdigtillverkade
      1 färdigutbildade
      2 färdigutvecklad
      1 färdigutvecklade
      1 färdigutvecklas
      1 färdigvuxen
      1 färdmedel
      1 färdriktningen
      1 färdvägar
      1 fåren
      2 fåret
      1 farfar
      2 farfara
     70 färg
      7 färga
      1 färgad
      8 färgade
      2 färgades
      3 färgämne
      9 färgämnen
      6 färgämnet
      1 färgändring
      4 färgar
     11 färgas
      3 färgat
      1 färgåtergivning
      1 färgats
      1 färgbilden
      1 färgblindhet
      1 färgdoppler
     40 färgen
     38 färger
      1 färgerna
      1 färgfällning
      1 färgförändringar
      1 färggranna
      1 färgkodad
      1 färgkodade
      1 färgkodning
      1 färgkontrasten
      1 färgkorrigeras
     17 färglös
     10 färglösa
      2 färglöst
      1 färgmättnaden
      1 färgmönster
      9 färgning
      1 färgningar
      1 färgningen
      1 färgningstekniken
      1 färgnyans
      3 färgpigment
      1 färgpigmenten
      1 färgpigmenter
      2 färgpigmentet
      1 färgsätta
      1 färgsätter
      3 färgseende
      1 färgskalans
      1 färgskiftningar
      1 färgskiftningen
      1 färgskrift
      2 färgstarka
      1 färgteckning
      1 färgtemperatur
      2 färgton
      1 färgvariationer
      1 färgytor
      1 farhågan
      4 farhågor
      1 farhågorna
      2 fårhund
      1 fårhundar
      1 farinae
      2 färjeläge
      1 fårklippare
      2 farkoster
     32 farlig
     39 farliga
      8 farligare
      1 farligast
      9 farligaste
      3 farlighet
      2 farligheten
     33 farligt
      4 farmaceuter
      3 farmaceutisk
      2 farmaceutiska
      4 farmaci
      2 farmacie
      1 farmacin
      1 farmaindustri
      3 farmaka
      2 farmakodynamik
      1 farmakodynamiken
      1 farmakodynamisk
      2 farmakodynamiska
      3 farmakokinetik
      1 farmakokinetiska
      1 farmakologer
     15 farmakologi
      1 farmakologikemi
      2 farmakologin
      1 farmakologins
     19 farmakologisk
      7 farmakologiska
      4 farmakologiskt
      4 farmakopé
      1 farmakopéen
      3 farmakopéer
      1 farmakopen
      7 farmakopén
      1 farmakoterapin
      5 farmakovigilans
      1 farmalogisk
      1 farmodern
      2 farmor
      1 färnebofjärden
      1 faroanalys
      8 faror
      6 fåror
      1 farozon
     37 färre
      1 fars
      7 färsk
      7 färska
      1 färskfryst
      1 färskmassa
      1 färskmassabaserade
      5 färskt
      1 färskvatten
      1 farsot
      4 farsoten
      1 farsoter
      1 farstukvisten
      1 fårstyng
     14 fart
      2 fårtarmar
      7 farten
      1 farthämmande
      6 farthinder
     15 fartyg
      1 fartygen
      4 fartyget
      1 farvatten
      1 faryngal
      2 faryngala
      4 faryngeal
      1 faryngeala
      6 faryngit
      2 farynx
     58 fas
     31 fås
      1 fasa
      1 fasadbeklädnad
      1 fasaden
      1 fasadens
      3 fasader
      1 fasats
      1 fasberoende
      4 fasceit
      1 fasci
      3 fascia
      1 fasciculata
      1 fasciculus
      1 fasciit
      1 fascikelblock
      1 fascination
      1 fascinerande
     30 fasen
     16 faser
      5 faserna
      1 fasförskjutning
      2 fasinformation
      1 fasinformationen
      1 fasläge
      1 fasoner
      1 fasor
      1 fass
      1 fasställas
      1 fasstudier
    121 fast
     11 fäst
     42 fasta
     22 fästa
      1 fästad
      1 fastade
      2 fastan
      8 fastän
      2 fästande
      1 fastans
      5 fastare
      7 fästas
      1 fastboende
     19 fäste
      1 fästeförlust
      1 fastemotorik
      2 fästen
      3 fästena
      1 fasteperioden
     29 fäster
      4 fästes
      1 fästet
      1 fastetid
      2 fastetiden
      1 fastfas
      1 fastigheten
      4 fastigheter
      1 fastighetsägaren
      1 fastighetsskötare
      1 fastighetsskötsel
      4 fästing
     11 fästingar
      3 fästingarna
      1 fästingart
      5 fästingbett
      1 fästingbettet
      5 fästingburen
      1 fästingburna
      4 fästingen
      2 fästingfeber
      1 fästinghalsband
      1 fästingpincett
      1 fastklämt
      2 fastlades
     11 fastna
      1 fastnade
     21 fastnar
      5 fastnat
      1 fästning
      1 fästpunkt
      1 fästpunkten
     15 fästs
      1 fastsätts
      3 fastslå
      1 fastslagit
      2 fastslagits
      4 fastslår
      1 fastslås
      7 fastslog
      1 fastslogs
      1 fastspänd
     27 fastställa
      5 fastställande
      1 fastställandet
      4 fastställas
      4 fastställd
      2 fastställdes
      3 fastställer
      6 fastställs
      4 fastställt
      6 fastställts
      1 fastväxning
      1 fästyta
      3 fat
     40 fåtal
      1 fatala
      1 fatale
      2 fåtaliga
      1 fate
      1 fatet
      1 fath
      7 fatigue
    172 fått
      5 fatta
      2 fattade
      1 fattades
      1 fattar
      2 fattas
      1 fattat
      2 fattig
     31 fattiga
      3 fattigare
      2 fattigaste
     10 fattigdom
      4 fattigdomen
      1 fattighus
      1 fattigläkare
      2 fattiglappar
      1 fattigsjukhus
      1 fattigt
      1 fatty
      1 fauchard
      1 faulks
      1 fauno
      1 faust
      1 faustparacelsus
      1 favoriserade
      1 favoritserie
      1 favoritsonen
      3 fbi
      1 fbis
      1 fcc
      1 fcrireceptorer
      1 fd
      1 f�d
     13 fda
      1 fdagodkänd
      1 fdas
      2 fdg
      4 fe
      1 feb
    187 feber
      1 feberattackerna
      1 feberbehandling
      1 feberfri
      3 feberfrossa
      1 feberinsjuknandet
      1 feberkramper
     17 febern
      6 febernedsättande
      1 febernedsättning
      1 febernvidare
      1 febernvirus
      3 febersjukdom
      2 feberstadiet
      1 feberstadium
      1 febertermometer
      1 febertoppar
      1 febervirus
      2 febr
      1 febris
     24 februari
      2 fecc
      2 feces
      1 federal
      3 federala
      3 federation
      1 federationen
      5 feedback
      1 feedbacksystem
      1 fehlings
      1 fejd
      3 fekal
      2 fekaloral
      1 fekalorala
      1 fekaltoralt
      1 fekundation
      1 fekunditet
     55 fel
     25 felaktig
     16 felaktiga
      3 felaktigheter
      1 felaktigheterna
     42 felaktigt
      1 felanvändande
      1 felbedömer
      1 felbehandlade
      1 felbehandlingar
      1 felden
      2 feldenkrais
      1 feldenkraismetoden
      1 feldenkreismetoden
      2 feldiagnoser
      1 feldiagnosticerats
      1 feldiagnosticeringar
      1 felen
      8 felet
      1 fellatio
      1 fellcin
      2 fellea
      3 felmarginal
      1 felmarginalen
      1 felmätta
      1 felplacerad
      1 felrapporterat
      1 felsätta
      1 felsökning
      2 felställda
      1 felställning
      3 felställningar
      1 felställningen
      1 felsväljning
      1 feltolkningar
      1 felvänd
      1 felvändbri
      1 felveckade
    156 fem
      1 femårig
      1 femårsöverlevnad
      5 femårsöverlevnaden
      1 femen
      1 femenaktioner
      1 femfaktorteorin
      1 femflikig
      2 femidom
      3 feminisation
      1 feminiserat
      1 feminismen
      1 feministen
      3 feminister
      1 feministiska
      1 femlingar
      1 femme
      1 femprocent
      1 femring
      1 femsex
      1 femtal
      1 femtaliga
     15 femte
      3 femtedel
      4 femtio
      1 femtiotal
      1 femtiotalet
      7 femton
      2 femtonde
      1 femtunga
      1 femtusen
      1 fenacetin
      1 fenan
      1 fenazopyridin
      2 fencyklidin
      1 fenestration
      1 fenestrerad
      2 fenestrerade
      1 fenetylamin
      1 fenetylamindroger
      1 fenetylaminer
      1 fenetylaminsläkting
      1 fengshui
      1 fenmetralin
      3 fenmetrazin
     18 fenol
      1 fenolatjonen
     11 fenoler
      1 fenolerna
      1 fenoleter
      1 fenolhbensotriazolylmetyl
      1 fenolsulfonsyra
      1 fenom
     55 fenomen
      2 fenomenen
     28 fenomenet
      1 fenomenets
      1 fenomenologin
      3 fenotyp
      1 fenotypdrag
      1 fenotypdragen
      2 fenotyper
      1 fenotyperna
      1 fenotypiska
      1 fentanyl
      2 fentiazinderivat
      1 fentolamin
      1 fen�tre
      1 fenylaceton
      1 fenylacetonet
      5 fenylalanin
      2 fenylalaninhydroxylas
      1 fenylalaninnivåer
      4 fenylalaninnivåerna
      1 fenylalkamin
      1 fenyletylamin
      1 fenyletylaminoketoner
      6 fenylketonuri
      2 fenylpropanolamin
      1 fenytoin
      2 feodala
      1 feofytin
      2 feokromocytom
      2 feomelanin
      4 ferdinand
      1 ferm
      1 fermentation
      1 fermenterad
      1 fermenterade
      2 fermenterar
      1 fermenteras
      8 fermentering
      2 fermenteringen
      1 fermenteringsprocessen
      5 feromon
     18 feromoner
      2 feromonerna
      2 feromoners
      2 feromonet
      1 ferranti
      1 ferrara
      1 ferrari
      1 ferredoxin
      4 ferritin
      1 ferritinkomplex
      1 ferritinmätningar
      1 ferrocyanider
      1 ferromagnesiumineraler
      2 ferrosan
      1 ferrosans
      1 ferroxidas
     19 fertil
     17 fertila
      1 fertilin
      1 fertilisera
      1 fertiliseras
      3 fertilisering
     21 fertilitet
      4 fertiliteten
      1 fertilitetens
      1 fertilitetsbehandlingar
      1 fertilitetsbehandlingarna
      1 fertilitetscykeln
      1 fertilitetskliniker
      1 fertilitetspåverkande
      1 fertilitetsproblem
      1 ferulifolia
      1 fesiooh
      1 festa
      1 festen
      1 festerna
      1 festivalen
      1 festligheterna
      1 festmåltider
      5 fet
     19 feta
      2 fetala
      2 fetalperioden
      5 fetalt
      3 fetare
      1 fethet
      1 fetisch
      1 fetischism
      1 fetischister
     99 fetma
      1 fetmaacceptansen
      1 fetmaepedemin
      4 fetmaepidemin
      1 fetmakontroversen
      8 fetman
      1 fetmans
      1 fetor
      1 fetstil
    104 fett
      1 fettämnen
      2 fettansamling
      1 fettbaserade
      3 fettbildning
      1 fettbildningen
      1 fettbubbla
      1 fettcellens
      5 fettceller
      5 fettcellerna
      1 fettdepå
      1 fettdistributionen
      3 fettdroppar
     19 fetter
      1 fetterfettliknande
      1 fetterna
     10 fettet
      4 fettets
      1 fettfärgning
      2 fettförbränning
      1 fetthaltig
      1 fetthinna
      2 fettinlagring
      2 fettinnehåll
      1 fettintag
      1 fettklumpar
      1 fettkonsumtionen
      1 fettlagrande
      2 fettlagret
      4 fettlever
      1 fettlöslig
     12 fettlösliga
      1 fettlöslighet
      1 fettlösligt
      1 fettmängd
      1 fettmetabolismen
      1 fettmolekyler
      2 fettnekros
      1 fettnivåer
      1 fettområdet
      1 fettoxidationen
      1 fettprodukter
      2 fettreserv
      1 fettreserven
      2 fettreserver
      1 fettrik
      1 fettrika
      2 fettsammansättning
      1 fettsnål
      1 fettsnåla
      1 fettsnålt
     13 fettsugning
      1 fettsugningen
      1 fettsvulst
      1 fettsyran
      2 fettsyrarester
      1 fettsyrasyntesen
      1 fettsyrekedjorna
     30 fettsyror
      1 fettsyrorna
      1 fettumörer
      1 fettupplösande
      3 fettväv
      3 fettväven
      9 fettvävnad
      1 fettvävnaden
      1 fettvävnader
      1 fettvävnaderna
      1 fettvävnanden
      1 fetu
      1 fetus
      1 feuchtersleben
      1 feuchterslebens
      5 fev
     10 fever
      1 fevvc
      3 ff
      3 ffa
      1 ffi
      1 ffrekvens
      5 fft
      1 fftalgoritmen
      1 fftanalysator
      1 ffv
      1 fg
      3 fgfr
      1 fgfrgenen
      2 fgv
      1 fh
      4 fiber
      1 fiberartade
      1 fibercementskivorna
      1 fiberdiametrar
      2 fiberendoskopisk
      2 fiberfattig
      1 fiberfyllda
      1 fiberintag
      3 fiberoptik
      1 fiberoptisk
      1 fiberoptiskt
      2 fiberrik
      2 fibertillskott
      1 fibrat
      1 fibrater
     18 fibrer
      6 fibrerna
      1 fibrernas
      1 fibriller
      1 fibrillerna
      1 fibrilt
     14 fibrin
      3 fibrinet
      2 fibrinets
      2 fibrinnät
     11 fibrinogen
      1 fibrinolys
      1 fibrinolysin
      1 fibrinolytiska
      1 fibrintrådar
      1 fibrintrådarna
      1 fibro
      1 fibroadenom
      2 fibroblast
      4 fibroblaster
      1 fibrohyalin
      1 fibroider
      3 fibrom
      7 fibromen
     21 fibromyalgi
      1 fibromyalgia
      1 fibromyalgipatienter
      1 fibromyalgismärtor
      1 fibromyalgisyndrom
      1 fibronectin
     26 fibros
      1 fibrös
      1 fibrosarkom
      1 fibrosbildning
      1 fibroser
      1 fibrosstadiet
      2 fibröst
      1 fibrotiserande
      1 fibrotisering
      1 fibrotiska
      1 fibularis
      2 ficino
    201 fick
      3 ficka
      2 fickan
      2 fickklaffarna
      1 ficklampa
      1 ficklampans
      1 fickmätningssond
      4 fickor
      1 fickorna
      1 ficosis
      1 fictionberättelser
      1 fictiongenren
      1 fictionkaraktär
      1 ficus
      1 field
      3 fiende
      2 fienden
      2 fiendens
     10 fiender
      1 fiendernas
      1 fientlig
      1 fientliga
      1 fientlighet
      3 fientligt
      1 fife
      1 fifes
      1 fifth
      2 fig
      1 fighting
      1 figo
      5 figur
      5 figuren
      5 figurer
      1 fikon
      2 fiktion
      2 fiktiv
      7 fiktiva
      1 fikusar
      1 fikussläktet
      1 fila
      2 filament
      1 filamentbildande
      1 filamenten
      2 filamentöst
      1 filantrop
      1 filantropisk
      2 filariasis
      1 filarioidea
      2 fildigitalis
      1 fildigitalisstorahultrumswedenjpgfingerborgsblomma
      2 filer
      2 filialapotek
      1 filiformes
      1 filiformis
      7 filippinerna
      1 filippus
      2 filler
      1 fillers
     27 film
      1 filmarkiv
      1 filmarkivet
      1 filmatiserats
      2 filmbildare
      1 filmbildaren
      1 filmbildning
     12 filmen
      1 filmens
     12 filmer
      1 filmerna
      1 filmindustri
      2 filmindustrin
      1 filminspelningar
      1 filmisk
      1 filmjölk
      1 filmning
      1 filmregissörer
      1 filmskapare
      1 filmstjärnan
      1 filmsymboliken
      1 filon
      8 filosofen
      2 filosofer
      1 filosoferande
     16 filosofi
      5 filosofin
      2 filosofisk
      6 filosofiska
      3 filosofiskt
      4 filoviridae
      3 filovirus
      1 filovirusets
      1 filreras
      1 filt
      1 filtar
     19 filter
      1 filterkategorier
      1 filterreningsgrader
      1 filtertyp
      1 filtertypen
      1 filtning
      1 filtrationsfunktion
      1 filtrationshastighet
      1 filtrationshastigheten
      2 filtren
      5 filtrera
      2 filtrerad
      1 filtrerade
      1 filtrerar
      5 filtreras
      9 filtrering
      1 filtreringsprocesser
      1 filtreringssteg
      1 filtreringstekniker
      1 filtrerpapper
      1 fimbrier
      1 fimea
      2 fimos
      2 fimosis
      5 fin
      4 fina
      1 finalen
      1 finanserna
      1 finansiell
      1 finansiera
      1 finansierad
      1 finansieras
      2 finansiering
      1 finansieringssätten
      7 finare
      3 finaste
      1 finesser
      2 finflikiga
      2 finfördelas
      1 finfördelat
      1 finfördelning
      1 fingar
      3 fingarette
     10 finger
      1 fingeravtryck
      1 fingerborg
      1 fingerborgsblomma
      1 fingerborgsblomman
      1 fingerborgslikande
      1 fingerborgsört
      1 fingerfärdighet
      1 fingerhatt
      1 fingerkroksdragning
      1 fingerlika
      1 fingernaglar
      1 fingernaglarna
      1 fingerneuronerna
      1 fingerskadorna
      1 fingersugning
      1 fingertapping
      1 fingertopp
      3 fingertoppar
      3 fingertopparna
      1 fingertoppen
      1 fingertryck
      1 fingervarmt
      3 fingervisning
     29 fingrar
     14 fingrarna
      2 fingrarnas
      1 fingrars
      1 fingrat
      1 fingren
      4 fingret
      1 fingretnär
      1 finhåriga
      5 finjustera
      1 finjustering
      1 finka
      1 finkänsligt
     65 finland
      4 finlands
      1 finländsk
      3 finländska
      1 finlandssvensk
      1 finlandssvenskan
      1 finlandssvenskasanitär
      2 finmotorik
      1 finmotoriken
      1 finn
     38 finna
      1 finnålsbiopsi
      3 finnar
      1 finnarakne
    119 finnas
      1 finnbygderna
     30 finner
      1 finnish
      1 finnmarken
   2173 finns
      1 finporig
      1 finporigt
      1 finprickiga
      9 finsk
     21 finska
      1 finskan
      1 finskans
      1 finskbesläktade
      1 finslipning
      8 fint
      1 fintrådig
      1 finurlig
      1 finurliga
      1 fioler
      2 firades
      1 firandet
      4 firas
      1 firats
      1 fire
      1 fireknappen
      1 firenzuoli
      3 firetumme
      1 firman
      1 firmanamnet
      4 firmicutes
      1 fis
      1 fischer
      1 fisher
      1 fishermans
     33 fisk
      1 fiskallergier
     23 fiskar
      1 fiskare
      1 fiskarna
      1 fiskarnas
      1 fiskarten
      1 fiskarter
      2 fiske
      1 fiskinsulin
      1 fiskolja
      1 fiskrens
      3 fissilt
      4 fission
      2 fissionera
      1 fissionfusionfission
      1 fissionladdning
      1 fissionsladdningar
      1 fissionsladningar
      1 fissionsprodukter
      1 fissionsvapen
      1 fissur
      1 fissurer
      1 fissurförsegla
      6 fistel
      1 fistelgång
      1 fistlar
      4 fitness
      1 fitzgerald
      1 fiveyearold
      2 fix
      4 fixa
      3 fixera
      1 fixerade
      5 fixeras
      7 fixering
      1 fixeringar
      1 fixeringarna
      1 fixeringen
      1 fixeringsplatta
      1 fjäder
      1 fjäderfä
      1 fjäderliknande
      1 fjädermyggornas
      3 fjädern
      1 fjädrande
      9 fjädrar
      2 fjädrarna
     13 fjäll
      2 fjälla
      1 fjällad
      4 fjällande
     11 fjällen
      3 fjällig
      1 fjällika
      3 fjällning
      1 fjällräv
      1 fjällskivling
      1 fjällskivlingar
      2 fjälltrakterna
      1 fjällvandring
      1 fjälster
     22 fjärde
     10 fjärdedel
      4 fjärdedelar
      1 fjärdhundra
      1 fjärilar
      1 fjärran
      1 fjärrblockering
      1 fjärrmetastas
      1 fjärrmetastaser
      2 fjärrpunkten
      1 fjärrskådande
      2 fjärrstyrda
      1 fjärt
      1 fjärvärmekulvertar
      1 fjättrad
      1 fjelebo
      1 fjolårsgräset
      2 fjorton
     64 fkr
      1 fkr�
      5 fl
      6 fläck
     23 fläckar
      5 fläckarna
      3 fläcken
      2 fläckfeber
      2 fläckiga
      7 fläcktyfus
      1 fläcktyfusepidemi
      2 fläckvis
      1 fläckvisa
      1 fläckvist
     10 fladdermöss
      1 fladdermössen
      1 fladdermus
      1 fladdermusart
      1 fladdermusarterna
      1 fladdrar
      8 fläder
      1 fläderbären
      1 fläderblomchampagne
      1 fläderblommorna
      1 fläderblomssaft
      1 flädern
      1 fläderns
      1 fläderskinn
      2 flagell
      1 flagellanterna
      1 flagellaten
      1 flagellens
      1 flageller
      1 flaggärt
      1 flaggärtssläktet
      1 flaggbränning
      1 flagna
      5 flagnar
      1 flagor
      1 fläkt
      4 fläktar
      1 fläktdöden
      1 fläkten
      1 fläktyta
      1 flamenco
      1 flamman
      2 flamskyddsmedel
      1 flamugnar
      2 flanell
      1 flanken
      3 flankerna
      1 flänsost
      1 flänspackningar
      1 flare
      2 flashbacks
      1 flaska
      7 flaskan
      1 flaskformad
      1 flaskhalsen
      1 fläskkött
      1 fläskläpp
      4 flaskor
      1 flaskorna
      3 flat
      1 flätade
      3 flatlöss
      2 flatlus
      5 flatlusen
      1 flatlusens
      1 flätor
      1 flatt
      5 flatulens
      1 flatulensen
      2 flatus
      1 flaviviridae
      3 flavivirus
      2 flavonoider
      1 flavovirens
      1 flaxa
      1 flebit
      2 flebografi
      1 fleckeri
      1 fleischmannia
      1 flektion
      2 fleming
      2 flemming
      1 flemmings
      1 flensost
    178 fler
    805 flera
      1 fleräggsmånglingar
     20 flerårig
      8 fleråriga
      2 flerbarnsbörd
      1 flerbarnsbörder
      2 flerbarnsfödsel
      2 flerbörd
      1 flerbördsdräktigheter
      1 flerbördsgraviditet
      5 flercelliga
      1 flerdimensionellt
      1 flerfamiljshus
      1 flerfunktionsnedsättning
      1 flergångsalternativ
      1 flergångsartikel
      2 flergångsartiklar
      1 flergångsbruk
      1 flergångsmenskoppar
      1 flergångsprodukter
      1 flerkanalsoscilloskop
      1 flerkomponentpåsar
      1 flerkomponentsystemet
      1 fleromättade
      2 fleromättat
      1 flerorgansvikt
      1 flerskiktade
      3 flerskiktat
     95 flertal
     37 flertalet
      3 flervärda
     15 flest
    435 flesta
      1 flewett
      1 flexi
      2 flexibel
      4 flexibelt
      1 flexibilatis
      7 flexibilitet
      4 flexibla
      1 flexiblare
      1 flexitarianer
      1 flexner
      3 flexura
      9 flicka
      9 flickan
      1 flicknamn
     44 flickor
      1 flickorkvinnor
      2 flickorna
      3 flickornas
      4 flickors
      1 flight
      1 flik
      1 flikade
      6 flikar
      1 flikarna
      1 flikarnas
      1 flikas
      3 flikiga
      1 flikigt
      5 flimmerhår
      2 flimmerhåren
      1 flimmerhårens
      1 flimmerhårsceller
      1 flimmerhårscellerna
      2 flimrande
      1 flimrar
      1 flingor
      1 flint
      1 flinta
      1 flintshire
      1 flit
      2 flitig
      3 flitiga
     15 flitigt
      1 flitpengen
      3 floaters
      1 floby
      2 floccosum
      2 flock
      1 flockades
      2 flockar
      3 flockblommiga
      1 flockelsläktet
      1 flocken
      1 flockimmunitet
      1 flocklar
      1 flocklika
      1 flockmedel
      1 flockulering
      1 flod
      4 flöda
      1 flödande
      4 flödar
      2 flodblindhet
     12 flöde
      2 floden
      3 flöden
      4 floder
      1 floderna
      5 flödescytometri
      2 flödescytometrin
      1 flödesglottogrammet
      2 flödeshastigheter
      1 flödeshinder
      1 flödesinformation
      1 flödeskurva
      1 flödesmätare
      1 flödesprofil
     17 flödet
      1 flödets
      1 flödevolym
      1 flodfåror
      1 flodin
      2 flög
      7 flora
      5 floran
      1 floras
      3 florens
      1 florentinskt
      1 florenzer
      2 florerar
      5 flores
      1 floresiensis
      1 florey
      4 florida
      1 floroglucinol
      2 flos
      1 flottans
      1 flottfläckar
      2 flottor
      2 flow
      1 flowmätare
      1 flucytosin
      1 fluency
      4 fluga
      5 flugan
      1 flugans
      3 flugfångare
      1 flugfångaren
      1 flugfri
      8 flugor
      4 flugorna
      1 flugornas
      1 flugseende
     10 flugsvamp
      2 flugsvampar
      3 fluid
      2 flukloxacillin
      1 flukonazol
      1 fluktuationer
      1 fluktuera
      1 flunitrazepam
     10 fluor
      1 fluorättiksyra
      1 fluorecence
      1 fluorescein
      1 fluoresceiner
      2 fluorescens
      1 fluorescensljuset
      2 fluorescent
      2 fluorescerande
      1 fluorid
      2 fluorklormetan
      1 fluorkoncentration
      1 fluorlack
      1 fluorlacka
      1 fluormängd
      1 fluornivån
      1 fluoroform
      3 fluorokinolon
      6 fluorokinoloner
      1 fluoroskopi
      2 fluorsköljning
      1 fluortriklormetan
      1 fluothane
      1 fluoviler
      2 fluoxetin
      1 flurbiprofen
      1 fluro
      1 flushing
      1 flutide
      5 fly
      3 flyg
      9 flyga
      1 flygaktivitet
      4 flygande
      2 flygbesprutning
      2 flygbolag
      1 flygbuller
      3 flyger
      2 flyget
      1 flygfält
      1 flygfobi
      1 flyghudar
      1 flygigt
      1 flygmedicinen
      3 flygning
      1 flygolyckor
     12 flygplan
      1 flygplanet
      1 flygplans
      1 flygplansolycka
      1 flygplatser
      1 flygresa
      4 flygresan
      3 flygresor
      1 flygtid
      1 flygtorn
      1 flygvärdinna
      1 flygverksamheten
      1 flying
      7 flykt
      5 flyktig
      5 flyktiga
      1 flyktigare
      1 flyktigheten
      2 flyktingar
      2 flynn
      3 flynneffekten
      1 flyr
      1 flyt
      1 flyta
     31 flytande
      6 flyter
      1 flytning
      9 flytningar
      1 flytningarna
      2 flytningen
      2 flytt
     13 flytta
      5 flyttade
      5 flyttades
     11 flyttar
      9 flyttas
      3 flyttat
      1 flyttbar
      1 flytträning
      1 flyttstäda
      1 flyttstädad
      3 flyttstädning
      1 fmband
      2 fmedelvärde
      1 fmls
      4 fmri
      1 fmristudie
      1 fms
      4 fn
     24 fnkonventionen
      1 fnläkare
      1 fnmedlemmar
      2 fnorganet
      1 fnorganisationer
      6 fnöske
      2 fnösket
      2 fnösktickan
      2 fnösktillverkning
     21 fns
      1 fnskylten
      1 fnsoldater
      1 fnvarianten
      1 foalswort
      1 foamcell
      1 foamcells
     68 fobi
      3 fobibehandling
      2 fobidiagnoser
     46 fobier
      1 fobierna
      1 fobiker
     10 fobin
      3 fobisk
      8 fobiska
      1 fobityper
      2 fobos
      1 fÖc
      1 focal
      2 focus
     78 föda
     40 födan
      1 födanbr
      7 födande
      3 födans
      9 födas
      9 född
     34 födda
      3 födde
      9 föddes
     11 födelse
      1 födelsebeviset
      1 födelsedag
      1 födelsedagar
      3 födelsedatum
      1 födelsekohort
      2 födelsemärke
      6 födelsemärken
      9 födelsen
      1 födelseögonblicket
      1 födelsestatistiken
      5 födelsetal
      4 födelsetalen
      4 födelsevikt
      1 födelsevikter
      3 foder
      6 föder
      6 foderblad
      3 foderbladen
      1 foderflikarnas
      1 foderlikt
      1 foderpipen
      1 foderplatser
      1 föderskor
      1 fodertuben
      1 fodervägran
      1 födoämen
      7 födoämne
     26 födoämnen
      1 födoämnesallergen
      9 födoämnesallergi
      3 födoämnesallergier
      2 födoämnesaversion
      5 födoämnesintolerans
     15 födoämnesöverkänslighet
      1 födoämnesreaktionen
      1 födoämnesreaktioner
      3 födoämnet
     10 födointag
      2 födointaget
      1 födokälla
      1 födomotiverat
      1 födosök
      1 fodral
      7 fodret
     52 föds
     13 födsel
     38 födseln
      1 födselvikt
      3 födslar
      3 fog
      3 föga
      6 fogar
      3 fogarna
      2 fogarnas
      2 fogdar
      1 fogen
      1 foglig
      1 fogliga
      4 foglossning
      3 foglossningen
      1 fogningar
      1 fohmfs
      1 fokal
      5 fokala
      1 fokaladhesioner
      1 fokalpunkt
      2 fokalpunkter
      1 fokalt
     38 fokus
      1 fokusen
     17 fokusera
      6 fokuserade
      3 fokuserades
     27 fokuserar
      3 fokuserat
      1 fokusering
      1 fokuseringspunkt
      1 folat
      1 foleykateter
      1 foliata
      1 folie
      2 folium
      1 följ
     38 följa
     17 följaktligen
    129 följande
      1 följanden
     15 följas
    245 följd
      2 följda
     16 följde
     15 följden
     14 följder
      8 följderna
      2 följdes
      1 följdlögn
     12 följdsjukdomar
      1 följdsymptom
      1 följdtillstånd
      1 följdverkningar
      1 följdverkningarna
     71 följer
     16 följs
      2 följsamhet
      2 följsamma
     30 följt
     38 folk
      1 folkbildning
      4 folkbokföring
      2 folkbokföringen
      1 folkdräkt
      1 folkdräkten
      1 folken
      1 folkens
      4 folket
      3 folkgrupper
     12 folkhälsa
      8 folkhälsan
      1 folkhälsoarbete
      4 folkhälsoarbetet
      1 folkhälsoåtgärder
      2 folkhälsoenkäten
      1 folkhälsoexperter
      1 folkhälsofrågor
      4 folkhälsoinstitut
      2 folkhälsoinstitutet
      2 folkhälsokommittén
      1 folkhälsoministrar
      4 folkhälsomyndigheten
      2 folkhälsomyndighetens
      1 folkhälsonivå
      1 folkhälsonutrition
      1 folkhälsoområdet
      1 folkhälsoplanerare
      3 folkhälsoproblem
      1 folkhälsoproblemen
      1 folkhälsoråd
      1 folkhälsorapporten
      1 folkhälsosamordnare
      1 folkhälsostrateg
      2 folkhälsovetenskap
      1 folkhälsovetenskapens
      2 folkhälsovetenskapliga
      1 folkkommunernas
      1 folklagren
      1 folklig
      5 folkliga
      1 folkligt
      2 folklore
      1 folkmängden
      1 folkmängdens
      3 folkmassor
      3 folkmedicin
      8 folkmedicinen
      4 folkmedicinens
      1 folkmediciner
      1 folkmedicinisk
      2 folkmedicinska
      1 folkminskningen
      1 folkmord
      1 folkmordet
      7 folkmun
      1 folkräkningen
      1 folkrepubliken
      1 folkrikaste
      1 folkrörelsetraditioni
      5 folks
      1 folksaga
      3 folksjukdom
      1 folksjukdomar
      1 folksjukdomarna
      1 folksjukdomen
      1 folkskaror
      1 folkskyggare
      2 folkslag
      1 folkslaget
      1 folkstammar
      1 folkstammen
      1 folkstorm
      1 folktandvård
      1 folktandvården
      4 folktro
      4 folktron
      1 folkuppfattning
      1 folkvandringstida
      7 föll
      1 follicular
      1 follikel
      1 follikelceller
      4 follikelcellerna
      1 follikelcysta
      1 follikelcystor
      3 follikeln
      9 follikelstimulerande
      1 follikeltillväxten
      5 folliklar
      1 folliklarna
      3 follikulär
      2 follikulit
      2 follikuliter
      1 föllings
      1 following
      9 folsyra
      1 folsyraantagonist
      1 folsyraberikades
      1 folsyrabrist
      1 folsyran
      3 folsyrasyntesen
      1 folsyreantagonist
      1 folsyreantagonister
      1 folsyresyntes
      2 fom
      1 fomepizol
      1 fomiter
      3 fonasteni
      9 fonation
      1 fonationen
      1 fonationsstyrka
      1 fond
      1 fondkommissioner
      3 fonem
      1 fonematiskt
      2 fonemen
      1 fonetik
      1 fonetisk
      5 fonetiska
      2 foniater
      1 foniaterÖnhläkare
      7 fonofobi
      1 fonofobikänslighet
      1 fonografiska
      1 fonologi
      2 fonologisk
      1 fonologiska
      2 fonologiskt
     12 fönster
      2 fönsterglas
      1 fönsterputs
      1 fönsterputsning
      1 fönstertittarsjuka
      4 fönstertittarsjukan
      1 fönstren
      9 fönstret
      2 fontanellen
      1 fontanellerna
      1 fontänhus
      2 fontänhusen
      1 fontänhuset
      1 fontänhusetfountain
     12 food
      1 foods
      2 foot
     30 for
   8683 för
     44 föra
      2 förädla
      2 förädlade
      1 förädlats
      3 förädling
      3 förakt
     12 förälder
     15 föräldern
      4 förälderns
      1 förälders
      2 föräldrabalken
      1 föräldrabunden
      1 föråldrad
      1 föråldrade
      1 föräldraföreningar
      1 föräldraförmågor
      2 föräldraförmågorna
      1 föräldrahem
      2 föräldrakompetens
      1 föräldraledighet
     60 föräldrar
      1 föräldrarcellerna
     35 föräldrarna
     11 föräldrarnas
      1 föräldraromvårdnadspersoners
      3 föräldrars
      1 föräldrarsomvårdnadspersoners
      1 föräldrarvårdare
      1 föräldrarvårdnadshavare
      3 föräldraskap
      1 föräldraskapet
      1 föräldraskattningar
      1 föräldrastil
      1 föräldrastöd
      1 föräldrastödsprogram
      1 föråldrat
      1 föräldraträning
      1 föräldraträningsprogram
      7 föräldrautbildning
      1 föräldrautbildningar
      3 föräldrautbildningarna
      2 föräldrautbildningsprogram
      1 föräldrautbildningsprogrammen
      1 förälska
      4 förälskad
      1 förälskelse
      2 foramen
      2 föränderliga
      1 föränderlighet
     28 förändra
     27 förändrad
     19 förändrade
      7 förändrades
     11 förändrar
     44 förändras
     19 förändrat
     14 förändrats
     54 förändring
    126 förändringar
     13 förändringarna
     12 förändringen
      1 förändringens
      1 förändringsförmåga
      1 förändringsförmågan
      1 förändringsprocessen
      1 förändringsprocesser
      1 förångare
      4 förångas
      1 föraningen
      1 förankra
      1 förankrad
      2 förankrade
      2 förankrar
      1 förankrat
      2 förankring
      4 föranleda
      4 föranledde
      6 föranleder
      1 föranleds
      4 föranlett
      1 föranstalta
      1 förärad
      1 föräras
      1 förarbete
     12 förare
      5 föraren
      1 förarens
      1 förares
      1 förarga
      1 förargelseväckande
      1 förarkabinhuvar
      1 förarsäten
     19 föras
      1 föratt
      8 förband
      2 förbandet
      1 förbandsduk
      1 förbandsplats
      2 förbandsplatsen
     58 förbättra
     19 förbättrad
     13 förbättrade
      3 förbättrades
     16 förbättrar
     29 förbättras
      8 förbättrat
      8 förbättrats
     18 förbättring
      9 förbättringar
      1 förbättringarna
      3 förbättringen
      1 förbättringsfasen
      1 förbehåll
      1 förbehållet
      1 förbehandlad
      1 förbenas
      4 förbereda
      2 förberedande
      1 förberedd
      2 förberedelse
      2 förberedelsen
      4 förberedelser
      1 förberedelserna
      3 förbereder
      1 förberedningar
      2 förbereds
      1 förbestämda
     11 förbi
      3 förbinda
      9 förbindelse
      2 förbindelsen
     10 förbindelser
      2 förbindelserna
      4 förbinder
      1 förbindning
      1 förbinds
      1 förbipasserande
      1 förbise
      1 förbisedd
      2 förbises
      1 förbisett
      3 förbjöd
     10 förbjöds
      5 förbjuda
      9 förbjuden
      4 förbjuder
     27 förbjudet
      1 förbjudit
      4 förbjudits
     10 förbjudna
      4 förbjuds
      7 förblev
      7 förbli
     16 förblir
      1 förblivit
      2 förblöder
      2 förblödning
      1 förbluffade
      4 förbränna
      1 förbränner
     13 förbränning
      3 förbränningen
      1 förbränningsanläggningar
      3 förbränningsmotor
      1 förbränningsmotorer
      1 förbränningsprocesser
      2 förbränns
      1 förbränt
      4 förbruka
      4 förbrukar
      3 förbrukas
      1 förbrukning
      3 förbrukningen
      1 förbrukningsartiklar
      3 förbrukningsdag
      1 förbrukningsdagen
      1 förbrukningsdelar
      1 förbrukningsmaterial
      1 förbrukningstid
      2 förbrukningsvaror
      1 förbrutit
      1 förbryllade
     36 förbud
      1 förbuden
      8 förbudet
      2 förbudsmärken
      1 förbudsorienterad
      1 förbudstro
      2 förbund
      6 förbunden
      7 förbundet
      1 förbundit
      3 förbundna
      1 förbunds
      1 förbundsavgiften
      1 förbygga
      2 förbyggande
      1 force
      1 forced
      2 forcera
      4 forcerad
      1 forcerade
      2 forcerat
      1 förda
      1 fördärv
      5 förde
      2 fördefinierade
     26 fördel
      4 fördela
      2 fördelad
      5 fördelade
      1 fördelades
      1 fördelaktig
      4 fördelaktiga
      1 fördelaktigast
      7 fördelaktigt
     28 fördelar
     13 fördelarna
      3 fördelas
     25 fördelen
      4 fördelning
      7 fördelningen
     10 fördes
      2 fördisponerad
      2 fördjupa
      4 fördjupade
      1 fördjupning
      1 fördjupningar
      1 fördold
      1 fördolda
      1 fordom
      1 fördöma
      4 fördomar
      2 fördömde
      1 fördömer
      1 fördomsfullhet
      1 fördömt
     20 fordon
      6 fordonet
      4 fordonsbränsle
      1 fordonsindustri
      1 fordra
      2 fordrade
      2 fordrades
      1 fördraget
      2 fordrar
     10 fordras
      1 fordringsägare
      1 fördriva
      1 fördrivas
      1 fördrivits
      5 fördröja
      3 fördröjas
      4 fördröjd
      4 fördröjda
      2 fördröjde
      3 fördröjning
      1 fördröjningstiden
      1 fördröjt
      2 fördubblades
      2 fördubblar
      2 fördubblats
      5 fördubbling
      2 fördubblingstid
      1 fordyces
      1 fördyrar
    166 före
      3 förebild
      1 förebildat
      2 förebilder
      2 förebråelser
      1 förebud
     66 förebygga
     97 förebyggande
     11 förebyggas
     12 förebygger
      1 förebyggnad
      1 förebyggning
      4 förebyggs
      1 förebyggt
      6 föredatum
      3 föredatumet
     15 föredra
      2 föredrag
      2 föredragna
     28 föredrar
      5 föredras
      1 föredrog
      1 föredrogs
      3 förefalla
     23 förefaller
      1 förefintlig
      3 föreföll
      1 föregå
     12 föregående
     14 föregångare
      1 föregångaren
      1 föregångarna
      2 föregångsman
      3 föregår
     14 föregås
      5 föregåtts
      1 föregick
      1 föregivna
      2 föregripa
      1 föregripande
      1 föregriper
      1 föregrips
     38 förekom
    118 förekomma
    143 förekommande
    615 förekommer
     37 förekommit
     97 förekomst
     86 förekomsten
      1 förekomster
      1 förekomsterna
      1 förelåg
      2 föreläsningar
      1 föreläste
     10 föreligga
      1 föreliggar
     54 föreligger
     79 föremål
      2 föremålen
      4 föremålet
      1 föremåls
      6 förena
      6 förenad
      9 förenade
      4 förenar
      7 förenas
      9 förenat
     53 förening
     34 föreningar
      1 föreningarna
     19 föreningen
      2 föreningens
      1 föreningsstället
      1 förenkl
      3 förenkla
      2 förenklad
      3 förenklade
     10 förenklat
      1 förenklats
      3 förenkling
      1 förenklingen
      2 förenlig
      1 förenliga
      4 förenligt
      2 forensisk
      9 förenta
      1 föreskifter
      1 föreskrev
      1 föreskrevs
      5 föreskrift
     23 föreskrifter
      3 föreskrifterna
      1 föreskrivas
      1 föreskriven
      2 föreskriver
      2 föreskrivet
      1 föreskrivit
      1 föreskrivits
      1 föreskrivna
      1 föreskrivning
      1 föreskrivs
      6 föreslå
      1 föreslagen
      9 föreslagit
     17 föreslagits
      5 föreslagna
     21 föreslår
      2 föreslås
     22 föreslog
      5 föreslogs
      2 förespråka
      3 förespråkade
      2 förespråkades
      7 förespråkar
     18 förespråkare
     14 förespråkarna
      1 förespråkat
      2 forest
      3 föreställande
      1 föreställde
      4 föreställer
      6 föreställning
     17 föreställningar
      4 föreställningarna
      1 föreställningen
      2 föreställningsförmåga
      1 föreställningslivet
      1 förestod
      1 förestods
      4 företa
     54 företag
     15 företagen
     34 företaget
      4 företagets
      1 företagsamhet
      1 företagsbot
      1 företagsekonomi
      1 företagsekonomiskt
      1 företagshälsovård
      1 företagsledare
      1 företagsnamnet
      1 företagsstyre
      1 företagsvision
      2 företar
      6 företas
      7 företeelse
      3 företeelsen
      6 företeelser
      1 företogs
      3 företräda
      6 företrädare
      1 företrädarna
      1 företrädd
      2 företräder
     23 företrädesvis
      1 företrätt
      1 föreutsättning
      3 förfader
      6 förfäder
      1 förfäderna
      1 förfäktade
      1 förfäktades
      1 förfäktar
      4 förfall
      1 förfallen
      1 förfallna
      1 förfalskad
      1 förfalskade
      1 förfalskningar
      1 förfalskningarna
      1 förfaranden
      3 förfarandet
      1 förfaraonernas
      2 förfas
      1 författande
     15 författare
     12 författaren
      2 författarens
      1 författarinan
      8 författarna
      1 författarnas
      2 författarskap
      2 författning
      3 författningar
      1 författningarna
      1 författningen
      1 författningsenligt
      3 författningssamling
      1 förfelat
      1 förfina
      1 förfinad
      2 förfinade
      1 förfinades
      1 förfinat
      1 förfinats
      3 förflutna
      1 förflyktigas
      2 förflyta
      2 förflyter
      9 förflytta
      1 förflyttande
      5 förflyttar
      6 förflyttas
      1 förflyttat
      1 förflyttats
      7 förflyttning
      4 förflyttningen
      1 förflyttningssätt
      1 förfogande
      1 förfogar
      5 förföljd
      1 förföljda
      1 förföljdes
      3 förföljelse
      1 förföljelseidéer
      2 förföljelsekänsla
      6 förföljelsemani
      2 förföljelser
      1 förföljelseupplevelse
      2 förföljer
      1 förför
      1 förförelseteori
      1 förförisk
      1 förförstärkare
      1 förfrusen
      2 förfrysning
      1 förfylld
      1 förgänglighet
      1 förgångna
      1 förgård
      1 förgasade
      1 förgasas
      1 förgasning
      1 forget
      8 förgifta
      2 förgiftad
      2 förgiftade
      2 förgiftades
      1 förgiftar
      3 förgiftas
      4 förgiftat
     64 förgiftning
     23 förgiftningar
      8 förgiftningen
      1 förgiftningöverdosering
      6 förgiftningsfall
      2 förgiftningsrisk
      1 förgiftningssymptomen
      2 förgiftningssymtom
      2 förgiftningstillståndet
      2 förgrenad
      2 förgrenade
      4 förgrenar
      1 förgrenas
      1 förgrening
      4 förgreningar
      1 förgreningspunkt
      1 förgripa
      1 förgrovning
      1 förgrundsgestalt
      1 förgrundsgestalter
      2 förgyllt
      3 förhålla
     54 förhållande
     53 förhållanden
     15 förhållandena
     23 förhållandet
     20 förhållandevis
      1 förhållandevisvanlig
      7 förhåller
      1 förhållningsregler
      7 förhållningssätt
      1 förhand
      2 förhandla
      1 förhandlingsuppgörelse
      1 förhandsbeställningar
      1 förhandstillstånd
      4 förhårdnad
      3 förhårdnade
      2 förhårdnader
      1 förhårdningar
      1 förhärskade
      2 förhärskande
      2 förhastat
      1 förhäxade
      1 förhäxat
    119 förhindra
      3 förhindrad
      3 förhindrade
      1 förhindrades
     38 förhindrar
     17 förhindras
      1 förhindrat
      1 förhindring
      1 förhistoria
      1 förhistorien
      4 förhistorisk
      2 förhistoriska
      1 förhöja
     63 förhöjd
     50 förhöjda
      2 förhöjning
     33 förhöjt
      2 förhoppning
      2 förhoppningar
      3 förhoppningen
      2 förhoppningsvis
      2 förhör
      1 förhöret
      1 förhorning
      1 förhörsmetoderna
      4 förhud
     30 förhuden
      2 förhudsförträngning
      1 förhudsplastik
      1 förindustriell
      1 förinställda
      1 förinställts
      1 förintade
      2 förintelseläger
      1 förintelsen
      1 förjagare
      1 förjäses
      1 förkalkade
      1 förkalkning
      1 förkämpe
      1 förkänningen
      1 förkasta
      3 förkastade
      2 förkastas
      1 förkastats
      1 förkastelse
      1 förkastlig
      1 förkastliga
      7 förkläde
      2 förkläden
      1 förklädet
      1 förklädets
     35 förklara
      8 förklarade
      2 förklarades
      1 förklarande
     19 förklarar
     32 förklaras
      4 förklarat
     41 förklaring
     17 förklaringar
      1 förklaringarna
     13 förklaringen
      6 förklaringsmodell
      2 förklaringsmodellen
      3 förklaringsmodeller
      1 förklaringssyfte
      2 förklarliga
      1 förknipat
      1 förknippa
     20 förknippad
     25 förknippade
      7 förknippades
     35 förknippas
     20 förknippat
      8 förknippats
      1 förkokning
      3 förkorta
      2 förkortad
      3 förkortade
      1 förkortades
      7 förkortar
      9 förkortas
     26 förkortat
     19 förkortning
      8 förkortningen
      3 förkristen
      2 förkroppsligade
      1 förkroppsligat
      1 förkrympt
      3 förkrympta
      1 förkunnare
      3 förkunskap
      1 förkunskaper
     54 förkylning
     16 förkylningar
      1 förkylningsrelaterad
      3 förkylningssymptom
      1 förkylningssymtom
      1 förkylningssymtomen
      4 förkylningsvirus
      1 förlades
      1 förlag
      1 förlåga
      1 förlagan
      1 förlagd
      1 förlagen
      1 förlägenhet
      1 förlaget
      1 förlägganden
      4 förlägger
      2 förläggs
      1 förlagt
      1 förlama
      2 förlamad
      4 förlamade
      3 förlamande
      1 förlamar
     24 förlamning
      8 förlamningar
      6 förlamningen
      1 förlamningssjukdom
      1 förlamningssjukdomar
      1 förlamningstillstånd
     10 förlänga
      1 förlängas
     10 förlängd
     18 förlängda
      3 förlänger
      4 förlängning
      1 förlängningar
      5 förlängningen
      1 förlängningsbehandlingar
      6 förlängs
      3 förlängt
      1 förlåtande
      1 förlåtna
      1 förled
      3 förleda
      2 förledet
      1 förlegade
      1 förligger
      1 förlika
      1 förliste
      2 förlita
      4 förlitar
      1 förlöjligande
      5 förlöpande
      2 förlöper
     31 förlopp
     13 förloppet
      1 förloppets
      1 förlöpte
     12 förlora
     14 förlorad
     18 förlorade
      1 förloradökad
     23 förlorar
      1 förloraren
      1 förlorarna
      4 förloras
     18 förlorat
      1 förlorats
      2 förlösas
     58 förlossning
     14 förlossningar
      3 förlossningarna
     62 förlossningen
      2 förlossningens
      2 förlossningsarbete
      1 förlossningsarbetet
      3 förlossningsavdelning
      1 förlossningsavdelningen
      1 förlossningsbiträde
      2 förlossningsdepression
      1 förlossningsinstrument
      1 förlossningskanalen
      1 förlossningskatastrofer
      1 förlossningsklinikerna
      1 förlossningskonstbarnmorskekonst
      2 förlossningskonsten
      2 förlossningsläkaren
      1 förlossningsliknande
      1 förlossningsmedicin
      2 förlossningsmetod
      1 förlossningsoperation
      1 förlossningsoperationerna
      1 förlossningsplanering
      1 förlossningspsykos
      1 förlossningspulver
      2 förlossningsrädda
      3 förlossningsrädsla
      1 förlossningsrummen
      2 förlossningsrummet
      1 förlossningssmärta
      1 förlossningstång
      1 förlossningstången
      1 förlossningstänger
      1 förlossningsvägen
      3 förlossningsvård
      4 förlossningsvården
      1 förlossningsväsende
      1 förlöst
      1 förlöste
      1 förlovning
     35 förlust
      9 förlusten
      2 förluster
    479 form
      7 forma
      4 förmå
      7 formad
      1 förmådde
      6 formade
    181 förmåga
    102 förmågan
      3 förmagarna
     17 förmågor
      3 förmågorna
     18 förmak
      9 förmaken
      3 förmakens
      1 förmaket
      1 förmaksdilatation
      1 förmaksfladder
      6 förmaksflimmer
      1 förmaksklaffarna
      1 förmaksstängningarna
     14 formaldehyd
      1 formaldehydsulfoxylsyra
      1 formalin
      1 formaliserade
      2 forman
     13 förmån
      3 formande
      1 formandet
      1 formändrande
      1 förmaningar
      7 formant
      1 formantbegrepp
      1 formanten
     10 formanter
      3 formanterna
      3 formanternas
      2 formantkaraktär
      1 formantkaraktären
      1 formantliknande
      1 formantsyntetiserare
      1 formantvärden
      8 formar
     15 förmår
      7 formas
      1 förmås
     13 format
      2 formatet
      2 formation
      9 formationen
      2 formationens
      1 förmått
      1 formbara
      1 formbart
      1 förmedeltid
      7 förmedla
      3 förmedlad
      2 förmedlade
      1 förmedlande
      9 förmedlar
      1 förmedlare
      5 förmedlas
      2 förmedlingen
      1 förmedlingscentral
      1 förmedveten
      5 förmedvetna
     11 formel
      1 formelenheter
     10 formell
      5 formella
      6 formellt
     45 formeln
    103 formen
    193 former
      1 formeringen
     23 formerna
      1 formgivna
      1 formgivningen
      2 förmildrande
      3 forminriktad
      1 förminska
      1 förminskad
      1 förminskade
      1 förminskas
      1 formlerna
      1 formliknande
      1 formning
      2 förmoda
      2 förmodad
      3 förmodade
      1 förmodan
      8 förmodas
      2 förmodat
      1 förmodats
      1 förmodern
      1 förmodliga
     21 förmodligen
      3 förmögenhet
      2 förmögna
      1 förmörkat
      1 formoterol
      1 formpressad
      2 formpressade
      1 formpressat
      1 formpressning
      1 formspråk
     19 formula
      1 formulakg
      1 formulär
      1 formuläret
      2 formulas
      1 formulation
      2 formulera
      5 formulerade
      3 formulerades
      1 formulerar
      1 formuleras
      2 formulerat
      3 formulering
      2 formuleringar
      1 formuleringarna
      1 formuleringen
      1 formuleringsåtgärder
      1 förmultnat
      1 formvariationen
      1 formyl
      3 förmyndare
      1 förmyndarskap
      1 förmyndarskapet
      1 förmyndarverksamhet
      1 förmynderskapsreform
      6 forna
      1 förnämligast
      1 förnamn
      1 förnärmade
      1 fornegyptiska
      1 förnekade
      2 förnekande
      6 förnekar
      1 förnekat
      1 förnekelse
      1 fornengelska
      3 fornfranska
      1 fornfranskans
      1 fornhögty
      3 förnimma
      2 förnimmas
      1 förnimmelsen
      3 förnimmelser
      1 forniriskans
      1 fornlågtyska
      2 fornnordisk
      2 fornnordiska
      1 fornnordiske
      5 fornsvenska
      1 fornsvenskan
      1 fornsvenskans
      4 forntida
      3 forntiden
      4 förnuft
      7 förnuftet
      2 förnuftig
      1 förnufts
      1 förnuftsmässigt
      1 förnya
      3 förnyad
      1 förnyade
      4 förnyas
      1 förnyat
      1 förnybar
      2 förnyelse
      5 förödande
     16 föröka
      2 förökad
     35 förökar
      3 förökas
     11 förökning
      3 förökningen
      1 förökningsmetod
      1 förolyckad
      1 förorättade
      1 förorda
      2 förordade
      2 förordades
      2 förordar
      1 förordas
      1 förordnades
      7 förordning
      2 förordningar
      4 förordningen
      3 förorenad
      6 förorenade
      1 förorenas
      6 förorenat
      1 förorenats
      4 förorening
     14 föroreningar
      1 föroreningarna
      8 förorsaka
      2 förorsakad
      3 förorsakade
      1 förorsakades
      1 förorsakande
     17 förorsakar
      4 förorsakas
      3 förorsakat
      3 förövaren
      2 förpackad
      1 förpackade
      1 förpackades
      1 förpackaren
      2 förpackas
      1 förpackat
      4 förpackning
      2 förpackningar
      1 förpackningarna
      5 förpackningen
      1 förpackningsdag
      1 förpackningsgas
      1 förpackningsprocedurerna
      1 förpassades
      1 förpliktigades
      1 förpraktik
      1 förprogrammerad
      1 förprogrammerade
      1 förpubertala
      1 förpuppa
      1 förpuppas
      1 förpuppning
      2 förpuppningen
     90 förr
     16 förra
      3 förråd
      1 förrädisk
      1 förrådsbefruktning
     60 förrän
      1 förrått
      1 förrättas
      1 forrnordiske
      1 förromersk
      1 förrullade
      5 förruttnelse
      1 förruttnelsen
      1 förruttnelseprocesser
     85 förs
      2 försåg
      4 försågs
      7 försäkra
      1 försäkrat
      1 försäkring
      2 försäkringar
      1 försäkringen
      1 försäkringens
      1 försäkringsbedrägerier
      2 försäkringsbolag
      2 försäkringsbolaget
      1 försäkringsbrevet
      9 försäkringskassan
      1 försäkringsliknande
      1 försäkringssystemet
      1 försäkringssystemets
      1 försäkringstagaren
      1 försäkringsutredningar
     16 försäljning
      1 försäljningar
     11 försäljningen
      2 försäljningsargument
      1 försäljningsökning
      1 försäljningsställen
      1 församling
      2 församlingen
      1 församlings
      8 försämra
     28 försämrad
      1 försämradförlorad
     14 försämrar
     20 försämras
      3 försämrat
      1 försämrats
     15 försämring
      2 försämringar
      3 försämringen
      1 försanthållen
      1 försatsen
      3 försatt
      2 försätta
      2 försättas
      6 försätter
      2 försätts
      1 forsberg
      7 förse
     19 försedd
     12 försedda
      1 försedimentering
      1 försedimenteringen
      2 förseglad
      1 förseglar
      1 försegling
      2 förseglingen
      4 försenad
      2 försenade
      1 försenades
      1 försenas
      1 försenat
      2 försening
      1 förseningen
      1 försensitiserat
     11 förser
      9 förses
      4 försett
      2 försetts
      8 försiktig
      3 försiktiga
     17 försiktighet
      1 försiktighetsåtgärd
      4 försiktighetsåtgärder
      2 försiktighetsmått
      5 försiktigt
      1 försjunkenhet
      1 försjunker
      4 forska
      2 forskade
      1 forskades
      1 förskämning
      4 forskar
      1 forskarbehörighet
      1 forskarbestämda
    102 forskare
     13 forskaren
      2 forskares
      1 forskargemenskapen
      6 forskargrupp
      3 forskargrupper
      2 forskarlaget
     24 forskarna
      1 forskarsjälen
      1 forskarskola
      1 forskarskolor
      3 forskarutbildning
      1 forskarutbildningar
      3 forskarvärlden
      6 forskas
      2 forskat
      3 forskats
      5 förskjuta
      1 förskjutbar
      2 förskjuten
      2 förskjuter
      1 förskjutet
      1 förskjutits
      3 förskjutning
      1 förskjutningen
      1 förskjuts
    224 forskning
      2 forskningar
      1 forskningdesto
     40 forskningen
      1 forskningens
      1 forsknings
      2 forskningsarbete
      1 forskningsartikel
      2 forskningsavdelning
      1 forskningsbaserat
      1 forskningschef
      1 forskningsdebatt
      4 forskningsevidens
      6 forskningsfält
      1 forskningsfynd
      2 forskningsgren
      1 forskningsingenjör
      1 forskningsinriktat
      1 forskningsinriktning
      1 forskningsinsatserna
      1 forskningsinstitutet
      1 forskningsintensiv
      1 forskningsintensivt
      1 forskningskemikalie
      2 forskningslaboratorier
      1 forskningslaboratorium
      1 forskningsläget
      1 forskningsmaterialet
      1 forskningsmedel
      2 forskningsmetoder
      1 forskningsmetoderna
      4 forskningsområde
      6 forskningsområden
      1 forskningsöversikt
      2 forskningsprojekt
      1 forskningsramprogram
      1 forskningsrapport
      1 forskningsreaktorer
      6 forskningsresultat
      2 forskningsresultaten
      1 forskningsresultatens
      1 forskningsrön
      1 forskningssammanhang
      2 forskningssammanställningar
      1 forskningsstöd
      1 forskningsstödet
      1 forskningsstudie
      1 forskningsstudier
      2 forskningssyften
      1 forskningsunderlag
      2 forskningsverksamhet
      2 förskola
      1 förskolan
      1 förskole
      3 förskoleåldern
      2 förskoleklass
      2 förskolepersonal
      2 förskolor
      2 försköna
      1 förskonat
      1 försköning
      1 förskrev
      4 förskriva
      3 förskrivas
      1 förskriven
      1 förskriver
      1 förskrivet
      1 förskrivna
      6 förskrivning
      1 förskrivningen
      1 förskrivningsorsaken
      2 förskrivningsrätt
      5 förskrivs
     15 förslag
      1 förslagen
      2 förslaget
      2 förslagsvis
      1 förslitning
      2 förslitningar
      3 förslitningsskada
      2 förslitningsskador
      1 försluta
      1 försluten
      1 försluter
      1 försöjer
     90 försök
     49 försöka
      1 försökdjurspersonal
      4 försöken
     85 försöker
     10 försöket
      1 försöks
      1 försöksbasis
     12 försöksdjur
      5 försöksdjuren
      1 försöksdjurens
      2 försöksgruppen
      1 försöksjournal
      1 försöksjur
      1 försöksobjekt
      1 försöksperson
      2 försökspersonen
      1 försökspersonens
      5 försökspersoner
      4 försökspersonerna
      2 försökspersonernas
      1 försöksprojekt
      2 försöksverksamhet
      1 försöksvis
     17 försökt
     21 försökte
      2 försommaren
      1 försorg
      3 försörja
      1 försörjas
      9 försörjer
      2 försörjningen
      2 försörjs
      1 förspänning
      1 förspillas
      1 förspråklig
      1 försprång
      2 forssell
      1 forsslund
    293 först
    744 första
     57 förstå
      1 förstabehandling
      1 förstådd
      4 förstådda
      1 förstadie
      5 förstadier
      1 förstadierna
      3 förstadiet
      9 förstadium
      1 förståeligt
     13 förståelse
      6 förståelsen
      1 förstående
      1 förstahandsalternativ
      3 förstahandsbehandling
      1 förstahandsbehandlingen
      1 förstahandsmedlen
      2 förstahandspreparat
      3 förstahandsval
      1 förstahandsvalet
      1 förstahjälpen
      1 förställningar
      1 förstämningsförändringar
      1 förstämningssyndrom
      2 förstånd
      1 förståndet
      3 förståndshandikapp
      2 förståndshandikappade
      1 förståndssvag
      1 förstapassagemetabolism
      2 förstapassagemetabolismen
      1 förstaplats
     11 förstår
     12 förstärka
      1 förstärkande
     11 förstärkare
      2 förstärkarens
      1 förstärkares
      2 förstärkas
      8 förstärker
     10 förstärkning
      1 förstärkningar
      1 förstärkningsfaktor
      7 förstärks
      8 förstärkt
      5 förstärkta
      1 förstärkte
     15 förstås
      1 förstaspråk
      1 förstatligad
      1 förstatligades
      1 förstavalsbehandlingen
     19 förste
      1 forsteri
      1 förstfödda
      1 förstfödde
      1 förstföderskor
      1 förstfödslorätten
      6 förstnämnda
      8 förstod
      1 förstods
      1 förstoppad
     21 förstoppning
     16 förstör
      6 förstora
      9 förstöra
     14 förstorad
     13 förstorade
      1 förstorades
      1 förstörande
      1 förstorar
      8 förstoras
      8 förstöras
      3 förstorat
      1 förstorats
      3 förstörd
      2 förstörda
      3 förstörelse
      4 förstoring
      2 förstoringar
      2 förstoringen
     22 förstörs
      4 förstört
      1 förstummas
      8 försumbar
      1 försumbart
      1 försumlig
      2 försumma
      2 försummade
      1 försummelsen
      3 försurning
      2 försvaga
      3 försvagad
      5 försvagade
      1 försvagades
      1 försvagande
      6 försvagar
      7 försvagas
     13 försvagat
      5 försvagats
      5 försvagning
      3 försvagningar
     11 försvann
     16 försvar
      8 försvara
      9 försvåra
      1 försvårad
      2 försvarar
     10 försvårar
      1 försvarare
      1 försvararna
      1 försvaras
      3 försvåras
      1 försvarat
      2 försvårat
      1 försvårats
      1 försvarbara
      6 försvaret
      1 forsvarets
      1 försvarsanläggningar
      1 försvarsbarriärer
      1 försvarsfunktionsskala
      1 försvarslinje
      1 försvarslösa
      3 försvarsmakten
      1 försvarsmaktens
      1 försvarsmek
      2 försvarsmekanism
      6 försvarsmekanismer
      1 försvarspolitik
      1 försvarsreaktion
      1 försvarsreaktioner
      1 försvarsrespons
      1 försvarsstaben
      1 försvarsstrategier
      2 försvarssystem
      1 försvarsystem
      1 försvenskats
     11 försvinna
     85 försvinner
      1 försvunna
      1 försvunnen
      1 försvunnet
     11 försvunnit
      1 forsyth
     36 fort
      1 for�t
      6 fört
      1 förtal
      1 förtär
      6 förtära
      1 förtärande
      6 förtäras
      1 förtärde
      2 förtärdes
     11 fortare
     21 förtäring
      4 förtärs
      2 förtärt
      1 förtärts
      1 förtas
      1 förtätning
      1 förtätningar
      2 fortbestånd
      1 fortbestår
      1 fortbilda
      1 fortbildningsnivå
     17 förteckning
      2 förteckningarna
      1 förteckningen
      1 fortfar
    166 fortfarande
      1 fortfor
      1 fortgå
      3 fortgående
      5 fortgår
      2 fortgick
     10 förtid
      2 förtida
      3 förtidig
      2 förtidsbörd
      1 förtidsbörden
      1 förtidspensionerade
      1 fortissimo
      1 förtjäna
      1 förtjänsttecken
      1 förtjänsttecknet
      4 förtjockad
      1 förtjockade
      1 förtjockare
      3 förtjockas
      3 förtjockning
      2 förtjockningar
      2 förtjockningen
      2 förtjockningsmedel
      1 fortledde
      3 fortlevnad
      1 fortlöpa
      5 fortlöpande
      2 fortlöper
      5 fortplanta
      1 fortplantade
      2 fortplantande
      7 fortplantar
      2 fortplantas
     30 fortplantning
      4 fortplantningen
      1 fortplantningenreproduktionen
      1 fortplantningsanpassningen
      1 fortplantningscykeln
      1 fortplantningsdriften
      1 fortplantningsförmåga
      1 fortplantningsförmågan
      4 fortplantningsorgan
      1 fortplantningsorganen
      1 fortplantningsorganens
      1 fortplantningssjukdomar
      7 fortplantningssystemet
      1 fortplantningssystemets
      2 förträfflighet
      1 förträgning
      2 förtränga
      1 förträngd
      2 förträngda
      8 förträngning
      4 förträngningar
      3 förträngningen
      3 förtroende
      2 förtroendet
      1 förtrollad
      2 förtrollningar
      8 förts
     31 fortsatt
      1 fortsätt
      9 fortsatta
     23 fortsätta
     15 fortsatte
      1 fortsätte
     43 fortsätter
      1 fortsattes
      3 fortsättning
      1 fortsättningar
      2 fortsättningen
      2 fortskred
      1 fortskrida
      5 fortskridande
      6 fortskrider
      1 fortskridit
      1 fortskridning
      1 fortstår
      1 förtunna
      1 förtunnats
      1 förtunning
      2 förtvålning
      1 förtvålningen
      1 förtvinade
      2 förtvinar
      4 förtvining
      1 förtvivlade
      2 förtvivlan
      2 förtydliga
      1 förtydligande
      8 forum
      1 forumen
      1 forumsida
      1 förunderligt
      1 förundersökning
      1 förundran
      2 förunnat
      6 förut
      2 förutbestämd
      2 förutbestämda
      1 förutbestämt
      2 förutfattade
      2 förutgående
    119 förutom
      3 förutsäga
      1 förutsägas
      3 förutsägbar
      1 förutsägbara
      1 förutsägbart
      1 förutsägelse
      1 förutsägelser
      1 förutsagt
      8 förutsatt
      1 förutsättande
      1 förutsättas
      1 förutsatte
     10 förutsätter
      1 förutsättes
     20 förutsättning
     32 förutsättningar
     11 förutsättningarna
      1 förutsättningen
      1 förutsatts
      2 förutse
      1 förutses
      2 förutspådde
      2 förutspås
      1 föruttnelse
      8 förväg
      1 förvägrats
      1 förvakuum
      1 förvällas
      2 förvällning
      1 förvaltar
      1 förvaltare
      1 förvaltas
      2 förvaltning
      1 förvaltningen
      1 förvaltningscykler
      1 förvaltningskunskap
      1 förvaltningskunskapen
      2 förvaltningslinje
      4 förvaltningslinjen
      2 förvaltningsmyndighet
      1 förvaltningsrätt
      1 förvaltningsuppgifter
      2 förvånade
      1 förvånades
      1 förvånande
      5 förvånansvärt
      1 förvandlad
      4 förvandlas
      2 förvandling
      1 förvåning
      1 förvanskad
      1 förvanskade
      2 förvanskning
      2 förvänta
      7 förväntad
      4 förväntade
      2 förväntades
      5 förväntan
      1 förväntar
     15 förväntas
      2 förväntat
      1 förväntbart
      1 förväntning
     11 förväntningar
      1 förväntningarna
      6 förvara
      1 förvarad
      1 förvarade
      1 förvarades
      1 förvarar
     25 förvaras
      2 förvarats
     11 förvaring
      1 förvaringsanvisningar
      1 förvaringsmetoder
      2 förvaringsplatsen
      1 förvaringstemperatur
      5 förvarning
     11 förvärra
      2 förvärrande
      9 förvärrar
     29 förvärras
      1 förvärrats
      7 förvärvad
     18 förvärvade
      1 förvärvande
      1 förvärvar
      1 förvärvas
      5 förvärvat
      4 förvärvats
      2 förvärvsarbetande
     10 förväxla
      1 förväxlar
     44 förväxlas
      1 förväxlat
      2 förväxlats
      1 förväxling
      1 förväxlingar
      1 förvedad
      1 förverkad
      1 förverkade
      3 förverkande
      1 förverkandeyrkande
      3 förverkliga
     11 förvildad
      3 förvildade
      2 förvildas
      1 förvillelserna
      3 förvirrad
      5 förvirrade
      1 förvirrande
      1 förvirrat
     24 förvirring
      1 förvirringen
      3 förvisso
      1 förvrängd
      1 förvrängda
      1 förvrängning
      1 förvrängningar
      2 förvriden
      1 föryngras
      2 föryngring
      1 föser
      4 fosfat
      1 fosfatas
      1 fosfatbrist
      1 fosfater
      1 fosfaterna
      3 fosfatgrupp
      1 fosfatgrupper
      1 fosfatgrupperna
      1 fosfatidylrest
      1 fosfatintoxikation
      1 fosfoglukomutas
      2 fosfokreatin
      1 fosfolipas
      1 fosfolipidbilagret
      6 fosfolipider
      1 fosfolipiderna
      1 fosfolipidlagret
      1 fosfoniumjodid
      1 fosfor
      1 fosforamidsenapsgas
      2 fosforescens
      1 fosforescerande
      1 fosformetabolism
      1 fosfors
      1 fosforskärmen
      1 fosforsyra
      1 fosforylasmutas
      1 fosforylera
      1 fosforylering
      1 fosforyleringar
      1 fosforyleringdefosforylering
      1 fosforyleringsmönstret
      1 fosforylkolin
      1 fosgen
      3 fossila
      1 fossilerna
     57 foster
      1 fosteranomali
      5 fosterdiagnostik
      2 fosterdiagnostiken
      3 fosterdöd
      2 fosterfett
      3 fosterfördrivande
      1 fosterhinnan
      1 fosterhinnor
      2 fosterhinnorna
      2 fosterhuvudet
      2 fosterlivet
      3 fosterperioden
      1 fosterrörelserna
      1 fosters
      1 fosterskada
      1 fosterskadande
      5 fosterskador
      1 fosterskadorna
     18 fosterstadiet
      1 fosterstadium
      1 fosterställning
      8 fostertiden
      6 fosterutveckling
     10 fosterutvecklingen
      4 fostervatten
      1 fostervattenden
      2 fostervattenprov
      1 fostervattensprov
      4 fostervattnet
      1 fostervecka
      1 fosterveckan
      2 fostra
      1 fostrade
      1 fostran
      1 fostre
      2 fostren
     62 fostret
     22 fostrets
      1 fóstri
     23 fot
      1 fotända
      1 fotbad
      1 fotbäddar
      1 fotboll
      1 fotbolls
      1 fotbollsarenorna
      1 fotbollsförbund
      1 fotbollsklubben
      2 fotbollsspelare
      1 fotbollsspelaren
      1 fotdiameter
     42 foten
     14 fotens
      2 fotfäste
      1 fothållning
      1 fothälsa
      1 fotisk
      1 fotkirurgi
      1 fotknölarna
      1 fotknölen
      2 fotleden
      1 fotledsrörelser
      1 fotliknande
      1 foto
      1 fotobiologin
      1 fotodetektor
      1 fotodimerisera
      1 fotoelektriska
      1 fotofilm
      2 fotofobi
      1 fotogenlyktor
      2 fotografera
      1 fotograferade
      1 fotografering
      1 fotografi
      2 fotografier
      1 fotografin
      1 fotografins
      6 fotografisk
      4 fotografiska
      2 fotografiskt
      1 fotografitekniken
      1 fotokatod
      1 fotokatoden
      1 fotokemiska
      1 fotokromiska
      1 fotolitografi
      1 fotolyseras
      2 fotomultiplikator
      1 fotomultiplikatorer
      1 fotomultiplikatorn
      1 fotomultiplikatorrör
      4 foton
      1 fotonenergi
      1 fotonenergier
      3 fotoner
      2 fotonerna
      1 fotoners
      2 fotonstrålning
      1 fotosensibilisering
      1 fotosensibilitet
      1 fotosyntes
      1 fotosyntesen
      1 fotosyntetiserande
      1 fototerapi
      1 fotpumpsdriven
      2 fotriktiga
      7 fotröta
      2 fotrötan
      1 fotryggen
      1 fots
      1 fotsår
      1 fotskena
      1 fotspåren
      4 fotsulan
      4 fotsulor
      9 fotsulorna
     13 fotsvamp
      1 fotsvampen
      1 fotsvapen
     16 fött
      1 fottåben
     27 fötter
     17 fötterna
      9 fötts
      1 fotvalv
      4 fotvalvet
      2 fotvalvets
      1 fotvalvsplattan
      1 fotvård
      2 fotvårtor
      1 fotzonterapi�reflexologiförbundet
      1 fou
      1 foucault
      1 fouenhet
      1 found
      9 foundation
      1 foundationbetald
      1 foundationpuder
      2 fountain
      2 fouriertransform
      1 fouriertransformanalysatorn
      1 fouriertransformation
      1 fouriertransformering
      1 fovea
      2 foveola
      1 fowleri
      5 fr
      1 fracastoro
      1 fracastoros
      1 frack
      2 fradga
      1 fradgande
      1 fraenkel
     69 fråga
      1 frågade
     37 frågan
      3 frågar
      1 frågebatterierna
      1 frågefeber
      6 frågeformulär
      2 frågeformuläret
      1 frågeområdena
      1 frågeställaren
      2 frågeställning
      1 frågeställningen
      1 fragile
      4 fragment
      2 fragmentala
      1 fragmenteras
      1 fragmentering
      1 fragmentet
      1 fragmin
     34 frågor
      4 frågorna
      1 fragrances
      1 fraiche
      6 fräknar
      1 fräknarna
      1 fräkne
      1 frakt
      2 frakta
      1 fraktalmönster
      1 fraktar
      2 fraktas
      3 fraktion
      1 fraktionen
      1 fraktioner
      5 fraktur
      1 frakturen
     12 frakturer
      1 frakturkirurgi
      1 frälsare
      1 frälsning
      2 frälst
    330 fram
      1 framända
     36 framåt
      1 framåtböjd
      1 framåtböjning
      1 framåtbuktande
      1 framåtvända
      3 frambenen
      1 frambesvärja
      5 framboesi
      1 framboise
      5 frambringa
      2 frambringar
      1 framework
      6 framfall
      3 framfart
      1 framföder
    217 framför
      2 framföra
    105 framförallt
      1 framföranden
      1 framförandes
      1 framföras
      1 framförda
      1 framförde
      1 framfördes
      2 framförs
      1 framfört
      8 framförts
      2 framförvarande
      1 framfötter
      1 framfötterna
      1 framfötts
     24 framgång
      6 framgångar
      1 framgången
      1 framgångsfaktorn
     12 framgångsrik
      9 framgångsrika
     16 framgångsrikt
      9 framgår
      1 framhålla
      6 framhåller
      2 framhållit
      2 framhållits
      1 framhålls
      1 framhärda
      1 framhärdande
      2 framhäva
      1 framhävdes
      2 framhäver
      1 framhävs
      1 framhjärnan
      1 framhjul
      2 framhöll
      1 framhölls
     18 främja
      2 främjande
      9 främjar
      1 främjas
      1 främjat
     31 framkalla
      6 framkallad
      4 framkallade
      2 framkallande
     14 framkallar
     16 framkallas
      1 framkallat
      1 framkallningsvätskor
      2 framkom
      1 framkomlig
      2 framkommer
      2 framkommit
      1 framkomsten
      2 framlade
      3 framlades
      1 framlagd
      1 framlägga
      2 framlägger
      1 främling
      2 främlingar
      1 främlingarna
      1 främlingars
      4 framlob
      3 frammana
      1 frammanar
      1 frammanat
     48 främmande
      1 främmandesituationen
      7 framme
      1 framodlade
      3 framöver
      1 framprovoceras
     25 främre
      1 framrusande
      5 framsida
      8 framsidan
      1 framsidans
      1 framsidor
      2 framskridande
      2 framskriden
      2 framskridet
      5 framskridna
    315 främst
     39 främsta
      6 framstående
     23 framställa
      1 framställan
      1 framställandet
     16 framställas
      5 framställd
      5 framställda
      6 framställde
     14 framställdes
      6 framställer
     72 framställning
      1 framställningar
      2 framställningen
      1 framställningsmetoden
      1 framställningsprocess
     41 framställs
      4 framställt
      6 framställts
      3 framstår
      2 främste
     16 framsteg
      1 framstegen
      1 framsticker
      2 framtagandet
      3 framtagen
      3 framtaget
      2 framtagna
      1 framtagning
      1 framtagningen
      2 framtänderna
      1 framtass
      5 framtid
     23 framtida
     16 framtiden
      1 framtidsfullmakt
      3 framtidstro
      7 framtill
      1 framtog
      2 framtogs
      5 framträda
     16 framträdande
      1 framträdandet
     12 framträder
      1 framtvingades
      1 framtvingas
      1 framväggsinfarkt
      1 framväxande
      5 framväxt
      2 framväxten
   2911 från
      3 frän
      3 fran�aise
      2 france
      1 francine
      4 francis
      1 francisco
      1 francisella
      1 franco
      1 frånfiltrerar
      1 frånfiltreras
      2 frångå
      1 frangula
      3 frank
      1 frankfurt
      1 franklin
      1 frånkopplad
     57 frankrike
      1 franksson
      1 frånluftskanaler
      2 frånluftstumlare
      1 fran�ois
      2 fran�oise
      1 franqueti
      1 frans
      1 fransesco
      1 frånsett
     12 fransk
     54 franska
      1 franskan
      8 franskans
      1 franskbelgiske
     11 franske
      1 franskindianska
      1 franskschweiziske
      1 franskschweiziskt
      1 fransksvenskt
      1 franskt
      1 fransktyska
      5 fransmannen
      1 fransson
      1 frånstötande
      1 frånstötning
      2 fransyskan
      1 fråntagen
      1 fråntagits
      1 fråntar
      1 fråntas
      1 fråntogs
      1 frantz
      4 frånvarande
     20 frånvaro
      2 frånvaron
      4 franz
      1 franzosen
      2 fras
      2 fräsch
      3 fräscha
      1 fräschare
      1 fräscht
      1 frasen
      6 fraser
      1 fräses
      8 frätande
      1 fräter
      1 frätskador
      4 fred
      1 fredagarna
      2 freddie
      1 frederic
      3 frederick
      1 fredlös
      2 fredrik
      1 fredriks
      1 fredsgatan
      1 fredsmärken
      1 fredspipor
      3 free
      1 freedom
      1 freeganism
      2 freeman
      2 frej
     41 frekvens
      1 frekvensband
      1 frekvensdomän
     18 frekvensen
     26 frekvenser
      2 frekvenserna
      1 frekvensgången
      1 frekvenskomponent
      2 frekvenskomponenter
      1 frekvensläge
      1 frekvensnoggrannhet
      1 frekvensomfång
      1 frekvensomfånget
      3 frekvensområde
      1 frekvensområdet
      4 frekvensräknare
      1 frekventa
      1 french
      6 frenulum
      3 freon
      1 fresenius
      1 frestelse
     41 freud
      2 freudiansk
      6 freudianska
      1 freudkritik
     15 freuds
     31 fri
     38 fria
      1 friade
      1 friare
      1 friargåvor
      3 fribas
      1 fribasen
      1 fribaser
      1 frid
      1 fridans
      1 fridlysningen
      4 fridlyst
      1 fridyker
      2 fridykning
      1 friedelcrafts
      1 friedländer
      1 friedländers
      1 friedlieb
      1 friedreichs
     15 friedrich
      1 friend
      1 friendly
      1 fries
      5 friganer
      1 friganerna
      1 friganernas
      2 friganism
      1 friganismen
      1 friganismens
      1 frige
      4 frigiditet
      1 frigjorda
      1 frigjorts
      7 frigör
      5 frigöra
      1 frigörande
      3 frigörandet
      2 frigöras
      2 frigörelse
      1 frigörelsens
     21 frigörs
      9 frihet
      1 friheten
      1 friheter
      1 frihetsälskare
      1 frihetsberövas
      1 friidrottare
      1 friidrottaren
      1 friidrottsanläggningar
      1 frikändes
      1 frikänner
      1 frikopplad
      1 frikopplare
      1 frikopplat
      1 frikostiga
      7 friktion
      4 friktionen
      1 friktionselement
      1 friktionsljud
      1 friktionsmaterial
      1 frilägga
      1 friläggs
      1 friland
      1 friluftsaktiviteter
      1 friluftsbad
      4 friluftsliv
      1 frimärken
      1 frimärkssamlare
      1 fris
      4 frisätta
      4 frisättas
     13 frisätter
     12 frisättning
      4 frisättningen
      1 frisättningshormon
      1 frisättningshormoner
      1 frisättningshormonet
      1 frisättningshormonkörtlarna
      1 frisatts
     32 frisätts
      1 frisimmande
     46 frisk
     94 friska
      7 friskare
      2 friskfaktorer
      1 friskförklarats
      1 friskförklaringen
      1 friskhälsosamt
      1 frisknat
     13 friskt
      4 friskvård
      1 friskvårdsarbete
      1 friskvårdseurytmi
      1 frisläppa
      1 frisläppande
      1 frisläppas
      1 frisläpper
      2 frisläppningen
      4 frisläpps
      1 frisläppta
      1 frisörer
      1 frispark
      1 fristad
      7 fristående
      1 friståendebänk
      1 fristilsskidåkning
      1 frisyrer
      1 fritaga
      1 fritera
      1 friterad
      2 frith
      7 fritid
      4 fritiden
      1 fritids
      3 fritidsaktiviteter
      1 fritidsbåtar
      1 fritidsbegreppet
      1 fritidsbostadsförsäkringar
      1 fritidsbullret
      1 fritidsfrågorna
      1 fritidskontor
      1 fritidsnämnd
      1 fritidssektorn
      1 fritidssnickerier
      1 fritidsträning
      1 fritillaria
     36 fritt
      1 frityrolja
      7 fritz
      1 fritzsche
      1 friuli
      1 frivårdsinspektör
      6 frivillig
      9 frivilliga
      1 frivillighet
      1 frivilligorganisationer
     10 frivilligt
      7 frö
      1 fröämnen
      1 fröbaljor
      1 frodades
      4 frodas
      1 fröderberg
      1 fröding
      1 fröer
      2 fröet
      1 fröets
      1 fröförökas
      1 fröhylle
      3 fröimplantation
      2 frökapseln
      1 frökapslarna
      1 fröken
      1 frolovii
      3 from
      1 frömjöl
      1 fromma
     21 frön
     18 fröna
      2 front
      1 frontal
      2 frontala
      1 frontalgyrus
      1 frontalis
      6 frontalloben
      1 frontallober
      3 frontalloberna
      2 frontallobsdemens
      1 frontalplan
      1 fronten
      1 frontier
      3 frontmatad
      1 frontotemporal
      1 frontotemporala
      1 frontsoldaters
      2 frösådd
      2 frösättning
     18 frossa
      1 frossare
      1 frossbrytningar
      1 frosseriet
      1 frost
      1 frostat
      1 frostbite
      1 frostegård
      1 frosteriskenius
      1 frostskada
      3 frostskador
      1 frostskyddsmedel
      2 frotté
      1 frottering
      1 fröväxter
      1 fröväxternas
      1 frövitan
      8 fru
      2 fruar
      2 frukost
      1 frukostflingor
     14 frukt
      3 fruktad
      5 fruktade
      2 fruktämne
      1 fruktämnen
      3 fruktämnet
      2 fruktan
      1 fruktanlagen
      1 fruktansvärd
      2 fruktansvärda
      1 fruktansvärt
      2 fruktar
      1 fruktaromer
      1 fruktbaljor
      1 fruktbara
      1 fruktbarhetsgud
      1 fruktbarhetsgudar
      1 fruktbarhetssymbol
      1 fruktbarhetssymboler
      1 fruktbart
      1 fruktblad
     22 frukten
     19 frukter
      1 frukterbär
      1 frukterianerna
      7 frukterna
      1 fruktfladdermöss
      1 fruktförband
      1 fruktifikativ
      2 fruktkärnor
      1 fruktköttet
      1 fruktkroppar
      4 fruktkropparna
      2 fruktkroppen
      2 fruktkroppens
      2 fruktodlingar
      1 fruktos
      1 fruktsaft
      2 fruktsamhet
      1 fruktsamheten
      1 fruktsamhetsproblem
      1 fruktsamhetstoppen
      1 fruktsamt
      1 fruktsmaker
      3 frun
      1 frus
      2 frusen
      2 frusenhet
      1 frustrerade
      1 fry
      2 frys
      3 frysa
      1 frysas
      1 frysbehandlas
      1 frysbehandling
      1 fryseffekt
      1 frysembryon
      1 frysen
      3 fryser
      2 fryses
      3 frysning
      1 frysningsapparat
      1 fryspunkt
      1 frysskyddsmedel
      1 fryssnitt
      5 fryst
      1 frysta
      1 frystorkning
      9 fsh
      1 f�stra
      1 ftaabs
      1 ftaleinfärgämnen
      1 ftld
      1 fuchsia
      1 fuchsinet
      3 fue
      1 fuel
      2 fujian
      1 fuksin
      8 fukt
      2 fukta
      3 fuktad
      1 fuktade
      2 fuktängar
      1 fuktare
      1 fuktaren
      3 fuktas
      1 fukten
      1 fuktförlust
      2 fuktgivande
     18 fuktig
     16 fuktiga
      3 fuktighet
      1 fuktighetsbalansen
      1 fuktighetsbevarande
      8 fuktigt
      1 fuktion
      1 fuktkammare
      2 fuktkräm
      3 fuktkrämer
      1 fuktning
      1 fuktsäkert
      1 fukushima
      1 ful
      3 fula
      1 fulbom
      3 fulhet
     33 full
      2 fulla
      1 fulladdat
      2 fulländning
      1 fullbad
      1 fullbildad
      5 fullbildade
      3 fullborda
      2 fullbordad
      3 fullbordade
      1 fullbordar
      2 fullbordas
      1 fullbordat
      1 fuller
      1 fullfjädrade
      7 fullfölja
      1 fullföljande
      1 fullföljer
      2 fullföljt
      1 fullföljts
      1 fullgågna
      1 fullgånget
      5 fullgångna
      2 fullgjort
      6 fullgod
      2 fullgoda
      1 fullgörande
      4 fullgott
      1 fullhudsbrännskada
      2 fullkomligt
      1 fullkornsbröd
      1 fullkornsprodukter
     12 fullmakt
      4 fullmakten
      2 fullmaktens
      2 fullmäktig
      1 fullmäktigen
      1 fullmaktsgivare
      4 fullmaktsgivaren
      2 fullmaktsgivarens
      1 fullmaktstagare
      4 fullmaktstagaren
      1 fullnarkos
      4 fullo
      1 fullödig
      1 fullödigt
      1 fullpackas
      1 fullseende
      1 fullskalig
      1 fullspektrumlysrör
     19 fullständig
      4 fullständiga
     26 fullständigt
     52 fullt
      1 fullvaccinerade
      1 fullvärdiga
      1 fullvärdigt
      3 fullvuxen
      6 fullvuxna
      2 fumaria
      1 fumariaarterna
      1 fumigatus
      1 fumlighet
      1 fumus
      1 functio
      1 functional
      1 fund
      4 fundamental
      1 fundamentala
      3 fundamentalt
      2 fundera
      3 funderar
      1 funderingar
      6 fundus
      1 funduskörtelpolyper
     72 fungera
     12 fungerade
     27 fungerande
    182 fungerar
      2 fungerat
      2 fungicid
      1 fungicider
      1 fungiformes
      1 funiculus
      1 funkar
    243 funktion
      1 funktionalismen
      5 funktionalitet
      1 funktionaliteten
     33 funktionell
     44 funktionella
      8 funktionellt
     34 funktionen
    103 funktioner
      8 funktionerna
      1 funktions
      1 funktionsättet
      1 funktionsbedömning
      2 funktionsbortfall
      1 funktionsdugligt
      2 funktionsförmåga
      2 funktionsgenerator
      2 funktionsgeneratorn
     13 funktionshinder
      6 funktionshindrade
      2 funktionshindrande
      1 funktionshindret
      1 funktionslös
      1 funktionsmaterial
      2 funktionsmedicin
      2 funktionsnedsatt
      3 funktionsnedsättande
     38 funktionsnedsättning
     27 funktionsnedsättningar
      2 funktionsnedsättningarna
      6 funktionsnedsättningen
      1 funktionsnivå
      1 funktionsprincipen
      3 funktionssäkerhet
      1 funktionssätt
      3 funktionsstörning
      2 funktionsstörningar
      1 funktionstestning
      1 funktionsundersökning
      1 funktionverkan
      7 funna
      1 funnen
      1 funnet
     26 funnit
     56 funnits
      2 für
      1 furan
      2 furanokumariner
      2 furanring
      1 furansidan
      2 furosemid
      1 furunculus
      3 furunkel
      1 furunkeln
      6 furunklar
      1 fusera
      4 fuserar
      1 fuseras
      2 fusidinsyra
      1 fusidinsyrakräm
      1 fusiforma
      1 fusiformis
      3 fusion
      1 fusionsladdningen
      1 fusionsvapen
     19 fusk
      1 fuskanteckning
      1 fuskare
      1 fusklapp
      1 fusklapparna
      1 fuskmetod
      1 fvckvoten
      1 fvp
      3 fvt
      1 fykobilin
      2 fylaxis
     11 fylla
      3 fyllas
      6 fylld
      9 fyllda
      1 fylldblommiga
      2 fyllde
      2 fylldes
      1 fyllekärringar
     18 fyller
      1 fyllig
      2 fylliga
      5 fylligare
      1 fylligt
      1 fyllmedel
      2 fyllnad
      1 fyllnaden
      1 fyllnadsmedel
      1 fyllnadstryck
      3 fyllning
      1 fyllningar
      1 fyllningsmaterial
     14 fylls
      9 fyllt
      1 fylogenetiska
      1 fyn
     30 fynd
      6 fynden
      3 fyndet
      1 fyndigheten
      1 fyndigheter
      1 fyndort
      1 fyndplatsen
      1 fynduppgift
      2 fynduppgiften
    191 fyra
      1 fyraårig
      1 fyrfotadjur
      1 fyrkant
      2 fyrkanten
      1 fyrkanter
      1 fyrkantig
      4 fyrkantiga
      1 fyrkantigt
      4 fyrkantvåg
      1 fyrlingar
      1 fyrpol
      1 fyrpolms
      1 fyrtalet
      1 fyrtaliga
      3 fyrtio
      1 fyrtiotal
      1 fyrtiotalistgenerationen
      1 fyrverkerier
      1 fyrverkerisatser
      8 fysik
      1 fysika
      5 fysikalisk
      9 fysikaliska
      1 fysikaliskkemiska
      1 fysikaliskt
      1 fysikeffekter
      4 fysiken
      1 fysiker
      4 fysikern
      1 fysikmotorer
      1 fysikprofessorn
      1 fysiologanalytiker
      1 fysiologen
      2 fysiologer
     34 fysiologi
      5 fysiologin
     17 fysiologisk
     36 fysiologiska
      1 fysiologiskhormonella
      8 fysiologiskt
      1 fysioplogi
      1 fysioterapi
    116 fysisk
    123 fysiska
      1 fysiskasociala
      1 fysiskpsykisk
     41 fysiskt
      2 fytoalexiner
      2 fytohormoner
      1 fytolsidokedjan
      5 fytoöstrogener
      2 fytoöstrogenrik
      1 fytoterapi
     36 g
      5 �g
    152 gå
      6 gaba
      1 gabaa
      4 gabareceptorer
      5 gabon
      1 gabor
      1 gadd
      1 gaddar
      1 gadden
      2 gadefeldt
      1 gadelius
      7 gående
      1 gage
      1 gagea
      2 gagna
      1 gagnar
      1 gagnat
      1 gagrupper
      1 galaktografi
      8 galaktorré
      1 galaktorrén
      5 galaktos
      5 galaktosemi
      1 galaktosfosfaturidyltransferas
      1 galaktosintaget
      1 galaktosintolerans
      2 galantamin
      1 galapagossköldpaddan
      1 gälar
      1 gälarna
      1 galaxen
      1 galbanum
      1 galderma
      6 galen
      1 galenisk
      1 galenochymica
      6 galenos
      3 galenskap
      2 galgar
      1 galge
      1 galgen
      2 gall
     30 galla
     19 gälla
      1 gallagul
      1 gallalkoholer
     18 gallan
     35 gällande
      1 gallans
      1 gallaslemblod
      1 gallbesvär
      3 gallblåsa
     33 gallblåsan
      2 gallblåsans
      4 gallblåsecancer
      2 gallblåsegången
     19 gällde
      1 galledaren
    226 gäller
      1 galleri
      1 galleriet
      1 gallerior
      2 gallery
      1 gallfärgämne
      1 gallfärgämnet
      1 gallfeber
      1 gallflödet
      1 gallgång
      8 gallgångarna
     15 gallgången
      2 gallgångens
      6 gallgångscancer
      2 gallgräs
      1 gallien
      1 gallinsufficiens
      1 galliske
      1 gallium
      2 gallo
      6 gallsalter
      5 gallstas
     10 gallsten
      4 gallstenar
      1 gallstenen
      1 gallstensdiagnos
      1 gallstensproblem
      5 gallsyra
      1 gallsyreupptag
      6 gallsyror
      3 gallsyrorna
      1 gallsyrornas
      3 gällt
      1 gallträdet
      2 galltvål
      1 gallussyra
      3 gallvägar
      2 gallvägarna
      6 galna
      1 galnebär
      1 gal�nochymica
      1 galoscher
      4 galt
      2 galton
      1 galtons
      1 galvaniserat
      1 galvanisering
      2 galvanisk
      1 galvanometer
      1 gamas
      1 gambia
      1 gambiense
      1 gamble
      1 gamblers
      3 gambling
      3 gambusia
      2 gamet
      1 gametangier
      8 gameter
      2 gameterna
      1 gameternas
      1 gametocyten
      1 gametocyterna
      1 gametofyt
      1 gametofyten
      1 gametofyter
      1 gametogenes
      1 gametogenesen
     95 gamla
      1 gamle
      1 gamles
      1 gamling
      1 gammaglobulin
      1 gammaglutamyltransferas
      2 gammainterferon
      2 gammakamera
      1 gammaknivsbestrålning
     51 gammal
      1 gammaldags
      1 gammalgrekiska
     13 gammalt
      1 gammaperiod
      4 gammastrålning
      1 gammavågor
      1 gamofyten
      1 gamofyter
      1 gamow
      1 gandhis
    131 gång
      1 gäng
      6 gångar
      3 gångarna
      1 gångegenskaper
    112 gången
      1 gångens
    163 gånger
      1 gångerdag
      1 gångerna
      1 ganges
      1 gånghjälpmedel
      1 gångjärn
      1 gångkläder
      1 ganglier
      4 ganglierna
      1 ganglion
      2 gångna
      1 gångprov
      2 gangrän
      1 gangränös
      1 gangrenösa
      1 gångrubbning
      6 gängse
      1 gångsträckan
      1 gångsträckor
      1 gångsvårigheter
      1 gångsystem
      1 gångväg
     91 ganska
      2 gapa
      2 gapet
    422 går
      1 garage
      1 garaget
      6 garantera
      1 garanterad
      4 garanterar
      2 garanterat
      2 garanti
      1 garantier
      1 garcía
      1 gard
      1 gård
      3 gårdar
      3 gardasil
      2 gården
      1 garderobsblomma
      2 garderobsblomman
      1 gardet
      1 gårdfarihandel
      5 gardiner
      4 gardner
      1 gärdsgårdsstör
      1 gareth
      1 garinii
      1 gariscochrane
     27 gärna
      1 garnhärva
      4 gärning
      5 gärningar
      1 gärningen
      1 gärningsman
      1 gärningsmän
      4 gärningsmannen
      2 gärningsmannens
      1 gärningstillfället
      1 garva
      1 garvämnen
      1 garvning
     38 gas
      1 gås
      1 gasade
      1 gasades
      1 gasar
      1 gasavgång
      2 gasbildande
      3 gasbildning
      1 gasbinda
      1 gasbindan
      2 gasblandningen
      1 gasblåsa
      1 gasblåsan
      4 gasblåsor
      1 gåsblod
      1 gasbrand
      4 gasbubblor
      2 gasbubblorna
      6 gasemboli
     21 gasen
      1 gasens
     22 gaser
      3 gaserna
      1 gasernas
      1 gasers
      2 gasfickor
      2 gasformen
      2 gasformigt
      2 gasfyllda
      5 gåshud
      1 gåshuden
      1 gasjoner
      8 gaskammare
      1 gaskamrarna
      1 gasmixturer
      6 gasning
      1 gäsp
      2 gäspa
      6 gäspar
      1 gaspare
      7 gasparutto
      3 gäspning
      3 gäspningar
      1 gäspningarna
      1 gäspningen
      1 gäspningsreflexen
      1 gasrikt
      1 gasspisar
      1 gassprängning
      1 gassvullen
      1 gastätat
      2 gåstativen
      2 gåstativet
      1 gästdialys
      2 gaster
      4 gäster
      1 gästerna
      1 gasters
      1 gästhandduk
      1 gastkramning
      1 gåstöd
      1 gastral
      1 gastrektomi
      2 gastric
      2 gästrikland
      1 gästriklands
      6 gastrin
      1 gastrinceller
      1 gastriner
      3 gastrit
      7 gastroenterit
      1 gastroenteriter
      1 gastroenterologer
      1 gastroenterologi
      1 gastroenterology
      2 gastroesofageal
      1 gastrointestinal
      2 gastrointestinala
      2 gastrointestinalt
      1 gastroknapp
      1 gastrokolisk
      3 gastrokoliska
      4 gastroskop
      4 gastroskopet
      9 gastroskopi
      3 gastroskopin
      1 gastrostomi
      1 gastrostomikateter
      1 gastrovaskulärhåla
      1 gastroviva
      1 gasugn
     10 gasutbyte
      8 gasutbytet
      1 gasutläckning
      1 gasvagn
      2 gasväv
      5 gata
      1 gåta
      4 gatan
      1 gates
      4 gator
      2 gatorna
     43 gått
      1 gatubilden
      1 gatupoliser
      2 gauge
      1 gaugetal
      1 gauntlet
      1 gauss
      1 gaussenheten
      1 gauthier
     79 gav
      1 gåva
      2 gävle
      1 gävleborgs
      2 gåvor
     26 gavs
      1 gay
      1 gaykultur
      1 gaylussac
      1 gaynor
      1 gazette
      1 gazi
      1 gb
      1 gbs
      1 gceller
     10 gcm
      2 gcs
      1 gdf
      1 gdl
      1 gdnf
    456 ge
      1 geber
      1 geckoödlor
      2 gedigen
      1 gediget
      2 gee
      3 geel
      2 gees
      1 geist
      1 gekiskans
      9 gel
      3 gelatin
      1 gelatinsilverplåtar
      2 gelé
      1 geléaktig
      2 geléartad
      1 gelébh
      1 geléfyllda
      1 gelékudden
      1 gelelektrofores
      1 geléliknande
      1 gelen
      5 geler
      1 geleringsmedel
      2 gelform
      2 gell
      1 gellius
      1 gelplugg
      1 gem
      1 gemen
      1 gemene
      1 gemener
     25 gemensam
      1 gemensamheter
     28 gemensamma
     51 gemensamt
      3 gemenskap
      1 gemenskapens
      1 gemenskaperna
      1 gemzell
     23 gen
      1 genans
      2 genant
      5 genast
      1 genchips
      1 gendarmeri
      1 gendarmerie
      3 gendarmeriets
      1 gendarmerikårer
      1 gendarmeriorganisation
      1 gendefekter
      2 gender
      1 gendermatoser
      4 gendiagnostik
      1 gene
     35 genen
      1 genens
     49 gener
      1 genera
      7 general
      3 generaldirektör
      1 generaldirektoratet
      1 generaldirektörens
      1 generalerna
      1 generalförsamling
      1 generalförsamlingarna
      1 generalförsamlingens
      1 generalisera
      3 generaliserad
      3 generaliserade
      1 generaliserande
      7 generaliserat
      1 generaliserbarhet
      3 generalisering
      1 generaliseringar
      1 generaliseringen
      1 generalistutbildning
      2 generalsekreterare
      1 generalspersoner
      1 generandi
      1 generar
      6 generation
      4 generationen
     12 generationens
      4 generationer
      2 generationstid
      2 generationsväxling
      1 generationsvirus
      1 generationsvis
      2 generator
      2 generatorer
     24 generell
     21 generella
     66 generellt
      9 generera
      1 genererandet
      9 genererar
     10 genereras
      3 genererat
      1 generika
      1 generiska
      8 generna
      1 geners
      2 genes
      2 genesis
     10 genetik
      2 genetiken
      1 genetikens
      1 genetikerna
     44 genetisk
     73 genetiska
     35 genetiskt
      1 genfaktor
      2 genfelet
      2 genförändringar
      1 genfragmentet
      1 genfrekvens
      3 gengäld
      3 geni
      1 génie
      2 genier
      2 geniet
      1 geniets
      1 genioglossus
      3 genital
      5 genitala
      2 genitalia
      1 genitaliautvecklingen
      1 genitalier
      2 genitalierna
      1 genitalt
      2 genitiv
      1 geniunt
      2 genius
      1 genkloning
      1 genkomplex
      2 genmaterial
      1 genmaterialet
      1 genmodifierade
      2 genmutation
      2 genmutationer
   2042 genom
      1 genomarbetade
      1 genomblödning
      1 genomborra
      2 genomborrar
      1 genomborrats
     13 genombrott
      6 genombrottet
      1 genomesam
      7 genomet
      1 genomfart
      1 genomflöde
      1 genomflytning
      7 genomför
     49 genomföra
      4 genomförande
      1 genomförandet
     25 genomföras
      1 genomförbar
      1 genomförbart
      7 genomförd
      6 genomförda
      7 genomförde
     13 genomfördes
     22 genomförs
      6 genomfört
      5 genomförts
     26 genomgå
      7 genomgående
      5 genomgång
      3 genomgångar
      5 genomgången
      2 genomgånget
     48 genomgår
     26 genomgått
     12 genomgick
      5 genomgripande
      1 genomlevas
      1 genomlevde
      1 genomlidit
      1 genomlopp
      1 genomlysningsbild
      1 genompasserande
      1 genomsågat
      1 genomskådar
      1 genomskärning
      1 genomskärs
      4 genomskinlig
      6 genomskinliga
      5 genomslag
      1 genomsläpplig
      4 genomsläppliga
     11 genomsläpplighet
      1 genomsläppligheten
      2 genomsläppligt
     33 genomsnitt
      3 genomsnittet
     11 genomsnittlig
     22 genomsnittliga
      3 genomsnittligt
      3 genomsnittsåldern
      1 genomsnittsbilen
      1 genomsnittsformel
      1 genomsnittsliga
      1 genomsnittstiden
      1 genomsöks
      1 genomstekas
      1 genomströmmas
      2 genomströmning
      1 genomtänkta
      1 genomtränga
      4 genomträngande
      1 genomtränglig
      1 genomträngning
      1 genotoxiska
      1 genotropin
      2 genotypen
      2 genotyper
      1 genparet
      1 genpool
      2 genpoolen
      2 genpooler
      2 genprodukt
      1 genre
      1 genreglering
      1 gens
      1 genskador
      2 gensvar
      1 genteknik
      1 gentekniken
     16 gentemot
      6 genterapi
      1 gentest
      1 gentlemannen
      1 gentranskription
      1 gentranskriptionen
      2 genu
      3 genua
      1 genuesarna
      1 genuesiska
      1 genuin
      1 genuina
      1 genuint
      4 genuppsättning
      1 genus
      6 genusmedicin
      1 genusmedicinskt
      3 genusperspektiv
      4 genuttryck
      1 genuttrycken
      1 genvariant
      2 genvarianter
      1 genvarianterna
      1 genvariationer
      3 gen�ve
      1 gen�vekonventionen
      2 gen�vekonventionerna
      1 geofysik
      1 geografer
      2 geografisk
      3 geografiska
      7 geografiskt
      1 geologin
      1 geologiska
      2 geometriska
      2 georg
      3 george
      1 georges
      1 georget
      3 georgia
      1 georgien
      1 georgii
      1 georgiska
      1 geotekniska
      1 geovetenskap
    652 ger
      1 gerald
      1 geraniol
      1 geranium
      1 geranylpyrofosfat
      1 gerard
      1 gerbil
      5 gerhard
      4 geriatrik
      1 geriatriken
      2 geriatriker
      1 geriatrikern
      1 geriatrikerns
      1 geriatrisk
      2 geriatriska
      1 gerillaodling
      1 gerillasoldater
      1 germ
      1 germansk
      3 germanska
      1 germicid
      3 germicida
      1 gernreich
      1 geron
      1 gerontolog
      6 gerontologi
      2 gerontologin
      1 gerontologiska
      1 gerontology
      2 gerry
      1 gersonmetoden
      1 gersons
    181 ges
      1 gesäll
      1 gesällprov
      1 geschichte
      1 gest
      3 gestagen
      2 gestagener
      1 gestageninjektion
      2 gestagentabletter
      5 gestalt
      1 gestalta
      3 gestaltakademin
      2 gestaltar
      2 gestaltas
      1 gestalten
      2 gestalter
      1 gestaltpsykologin
      1 gestaltref
      3 gestaltterapeuter
      1 gestaltterapeutiska
      1 gestaltterapeututbildningen
      2 gestaltterapi
     14 gestaltterapin
      1 gestaltterapins
      1 gestationsåldern
      1 gestationsdiabetes
      3 gester
      5 get
      1 getah
      1 geten
      2 geting
      1 getingallergi
      7 getingar
      1 getingarbr
      1 getingen
      1 getinggift
      2 getingstick
      1 getingsting
      1 getmjölk
      1 getpors
      1 getrams
      1 gets
      1 getskinnskalsong
     30 gett
      5 getter
      2 getts
      1 geusis
      2 gevär
      1 gevärskulor
      5 gévaudan
      1 gévaudanmonstret
      3 gezondheidsraad
      2 gfaktor
      1 gfr
      1 ggc
      2 ggr
      1 ggt
      4 gh
      1 ghadenom
      1 ghana
      1 ghanaunder
      1 ghb
      1 ghee
      1 ghonfokus
      1 ghp
      2 ghrelin
      1 ghrh
      1 ghutsöndring
      2 ghz
      1 gi
      1 giant
      1 giardia
      2 giardiasis
      1 gibb
      1 gibberelliner
      1 gibboner
      1 gicht
     64 gick
      2 gid
      1 giddens
      1 giemsafärgning
     64 gift
      7 gifta
      1 giftärtor
      1 giftbägare
      1 giftbägaren
      1 giftblad
      2 giftblåsa
      1 giftchampinjon
      1 giftdos
      2 gifte
      1 gifteffekt
      1 gifteffekten
     39 gifter
      7 giftermål
      1 giftermålen
      1 giftermålet
      7 gifterna
     31 giftet
      1 giftfri
      2 giftfria
     64 giftig
     64 giftiga
      5 giftigare
      1 giftigast
      3 giftigaste
     19 giftighet
      4 giftigheten
      1 giftighetsgrad
     33 giftigt
      1 giftinformation
      1 giftinformationscentral
      7 giftinformationscentralen
     10 giftinjektion
      1 giftinjektioner
      1 giftkörtlar
      1 giftkörtlarna
      3 giftkremla
      2 giftkremlan
      1 giftmord
      1 giftmördad
      1 giftödla
      1 giftödlor
      1 giftorm
      1 giftproducerande
      1 giftproduktionen
      1 giftsnok
      2 giftsnokar
      1 giftstadgan
     21 giftstruma
      4 giftsumak
      1 giftsvamp
      1 giftsvamparna
     10 giftverkan
      1 giga
      2 giganteum
      3 giganteus
      2 gigantiska
      8 gigantism
      8 gigantomasti
      3 gigantomastin
      1 gigartina
      1 gikanalen
      1 gikanalens
     25 gikt
      1 giktbehandling
      1 gikten
      1 gilamonster
      1 gilaödla
      6 gilaödlan
      1 gilberts
      2 gilford
      2 gilgamesheposet
      4 gili
      1 giljotin
      1 gilla
      2 gillar
      1 gillas
      5 gillberg
      1 gillen
      1 gillette
      2 giltig
      2 giltiga
      2 gimetoden
      1 ginetex
      9 gingivit
      1 gingiviter
      3 ginkgo
      1 ginkgoÄven
      1 giona
      1 giovanni
      4 gips
      1 gipsbandage
      1 gipsningarna
      1 giriga
      1 girighet
      1 girl
      1 girls
      2 girolamo
      1 gissar
      4 gissel
      2 gisslan
      1 gisslande
     11 gisslarna
      1 gisslarnas
      2 gisslartågen
      1 gisslartåget
      1 gisslet
      1 gissning
      1 gissningar
      1 gissningsläser
      1 gitarrbyggaren
      1 gitarren
      1 gitarrens
      1 gitarrer
      1 gitarrist
      2 githago
      1 giva
      2 givande
      1 givärde
      5 givare
      1 givares
      1 givarland
      1 givarländer
      1 givarområde
      1 givarsystem
      5 given
     11 givet
      3 givetvis
     16 givit
      5 givits
      1 givmild
      4 givna
     37 gjord
     23 gjorda
     98 gjorde
     48 gjordes
     71 gjort
     36 gjorts
      1 gjörwellsgatan
      1 gjuta
      1 gjutas
      2 gjutjärn
      1 gjutna
      1 gjutning
      1 gjutningen
      2 gjuts
      1 gkg
      1 gkryptor
      1 �gl
      1 glaber
      2 glaciär
      1 glaciärolyckor
      2 glad
      1 glada
      2 gladare
      1 gladiatorer
      1 gladiatorerna
      1 glädja
      7 glädje
      1 glädjelöshet
      1 gladman
      2 gland
      2 glandel
      1 glandispapler
      2 glandler
      3 glandula
      2 glandulae
      1 glandulär
      1 glandulära
      4 glans
     10 glänsande
      3 glansig
      1 glansiga
      1 glansigare
      1 glansstrimmor
      1 glap
      1 glareolus
     72 glas
      1 glasbägare
      1 glasbjörk
      7 glasen
     19 glaset
      1 glasfibrer
      1 glasflaskans
      2 glasflaskor
      1 glasfönster
      1 glasföregångare
      6 glasgow
      1 glasgows
      1 glasgowskalan
      1 glasinfattningar
      1 glasinfattningarna
      2 glaskärl
      1 glaskonstnär
      5 glaskroppen
      3 glaskroppsavlossning
      1 glaskroppsavlossningar
      1 glaskroppsavlossningen
      1 glasmaterial
     31 glasögon
      5 glasögonbågar
      1 glasögonbåge
      1 glasögonbärare
      6 glasögonen
      1 glasögonframställningen
      2 glasögonglas
      1 glasögonmodet
      1 glasögonskalmar
      1 glasögontypen
      1 glasomvandlingstemperaturen
      1 glasoptik
      1 glasplåt
      6 glasplåtar
      2 glasplåtarna
      2 glasplåten
      1 glasrör
      1 glasruta
      4 glass
      1 glassfabriker
      1 glassföretag
      1 glassföretaget
      1 glassindustrin
      1 glasskiva
      1 glasskivor
      1 glassmärke
      1 glassmärken
      1 glasstillverkare
     11 glatt
      8 glatta
      1 glätta
      2 glättestenar
      1 glättning
      2 glättstenar
      2 glaubersalt
      7 glaukom
      1 glaukomformen
      1 glaukomsjukdomen
      4 glaxosmithkline
      1 glechoma
      1 glenn
      3 glesa
      1 glesare
      1 glesbygd
      1 glesbygdsmedicin
      3 glest
      1 gliacell
      3 gliaceller
      4 gliadin
      1 gliadinantikroppar
      1 gliadiner
      1 glida
      1 glidande
      2 glidat
      7 glider
      6 glidmedel
      1 glimmar
      1 glimsläktet
      2 glioblastom
      1 gliom
      1 glios
      1 glipar
      1 glis
      1 glitter
     17 global
      9 globala
      1 globalisering
     31 globalt
      1 globen
      3 globin
      1 �globin
      2 globinet
      1 globulärt
      9 globulin
      1 globulinvärden
      1 glock
      2 glöda
      3 glödande
      1 glödgning
      1 glödgningsresterna
      1 glödkatod
      2 glödlampor
      1 glödnät
      2 glödtråden
      2 gloeilampenfabrieken
      1 gloeospermus
      1 glomangiosarkom
      1 glömd
      1 glömde
      1 glömdes
      1 glomerulär
      1 glomerulära
      5 glomeruli
      3 glomerulonefrit
      1 glomerulonefriten
      1 glomerulosa
      1 glomeruloskleros
      1 glomerulus
      4 glömma
      4 glömmer
      1 glömsk
      3 glömska
      5 glömt
      1 glorifierar
      1 glorifieringar
      2 glossina
      2 glossit
      1 glossiten
      1 glossofobi
      1 glossopharyngealnerven
      1 glottidis
      4 glottis
      1 glottisöppning
      1 glottisstängning
      1 glottisvibrationerna
      1 gloucester
      1 glucose
      1 glue
      3 gluggar
     20 glukagon
      4 glukagonet
      1 glukagonets
      1 glukagonspruta
      1 glukan
      6 glukokortikoider
      1 glukokortikoidreceptorer
      5 glukoneogenes
      5 glukoneogenesen
      2 glukonsyra
     80 glukos
      2 �glukos
      1 glukosbrist
      2 glukosen
      1 glukosenhet
      1 glukosenheterna
      1 glukoset
      8 glukosfosfat
      1 glukosfosfatmolekylen
      1 glukosgalaktosmalabsorption
      1 glukoshalten
      1 glukoshalter
      1 glukosintolerans
      2 glukoskoncentration
      2 glukoskoncentrationen
      1 glukoskontroll
      3 glukosmätning
      1 glukosmolekyl
      1 glukosmolekylens
      2 glukosmolekyler
      1 glukosmonomerer
      1 glukosnivå
      1 glukosnivåer
      2 glukosnivåerna
      2 glukosnivån
      1 glukosreserven
      1 glukosrik
      1 glukossirap
      1 glukosvärdena
      1 glukuronater
      1 glukuronatjon
      3 glukuronsyra
      2 glut
      6 glutamat
      1 glutamatdehydrogenas
      1 glutamatinbindning
      1 glutamatkoncentrationen
      1 glutamatreceptorerna
      1 glutamatsemialdehyd
      2 glutamin
      1 glutaminas
      1 glutaminerg
      1 glutaminerga
      3 glutaminsyra
      1 glutamyltrna
      1 glutein
      1 gluteintolerans
     12 gluten
      1 glutenallergi
      1 glutenantikroppar
      1 glutenfri
      5 glutenfria
      2 glutenfritt
     15 glutenintolerans
      1 glutenintoleransen
      2 glutenintolerant
      2 glutenintoleranta
      1 gluteusmuskulaturen
      1 glycemiskt
      8 glycerin
      1 glycerinextrakt
     12 glycerol
      1 glyceroldel
      2 glyceroltrierukat
      1 glyceroltrioleat
      2 glyceryl
      1 glycerylstearat
      1 glycin
      1 glycinets
      2 glyfosat
      1 glyfosatbaserat
      1 glyfosyfat
      2 glykemiskt
     25 glykogen
      1 glykogenesen
      3 glykogenfosforylas
      1 glykogenfosforylaset
      1 glykogenin
      1 glykogennedbrytningen
      3 glykogenolys
      1 glykogenolysen
      1 glykogenreglerande
      3 glykogensyntas
      1 glykogensyntaset
      1 glykogensyntesen
      6 glykol
      1 glykolaldehyd
      1 glykoler
      1 glykolförgiftning
      1 glykolsyra
      1 glykolvin
      4 glykolys
      3 glykolysen
      1 glykolytiska
      6 glykopeptider
      1 glykopeptidresistens
      1 glykopeptier
      7 glykoprotein
      9 glykoproteiner
      1 glykoproteinerna
      1 glykoproteinet
      1 glykoproteinhormon
      1 glykoproteinkomplex
      1 glykoproteinlager
      1 glykoproteinreceptor
      3 glykos
      3 glykosid
      1 �glykosidbindingar
      3 glykosider
      1 gmelinii
      2 gmol
      4 gmr
      3 gmvolym
      1 gmvolymen
     24 gnagare
      2 gnagaren
      1 gnagarens
      1 gnagares
      1 gnager
      1 gnathostoma
      1 gned
      1 gnet
      2 gnetophyta
      1 gnetter
      4 gnida
      1 gnidas
      3 gnider
      2 gnidning
      1 gnidningar
      1 gnidningsljud
      1 gnidningsljudet
      3 gnids
      1 gnidstenar
      2 gnisslar
      1 gnisslare
      1 gnissling
      1 gnistbildande
      1 gnōmon
      1 gnosis
      5 gnrh
      1 gnrhanaloger
      4 gnugga
      1 gnuggande
      2 gnuggar
      2 gnyende
      1 goalball
    115 god
     55 goda
      1 göda
      1 godare
     17 godartad
     16 godartade
      2 godartat
      1 godartde
      1 godas
      1 gödas
      1 godenholm
      1 godfrey
      1 godhet
      1 godheten
      3 godis
      1 godiskonsumtion
     21 godkänd
     18 godkända
      1 godkände
      7 godkändes
      1 godkänna
      8 godkännande
      1 godkännanden
      4 godkännas
      2 godkänner
      2 godkänns
     12 godkänt
      7 godkänts
      1 gödning
      1 gödningsmedel
      1 godronii
      1 gods
      1 godsägare
      1 godsägarna
      2 gödsel
      7 godset
      1 gödsla
      2 godt
      1 godtagbara
      4 godtagbart
      1 godtroende
      1 godtrogen
      1 godtycke
      2 godtycklig
      1 godtycklighet
      1 godtyckligt
      2 godwin
      1 goes
      2 goethe
      1 goethes
      1 gogh
      1 goiter
      1 goitrogener
      1 gökärt
      1 gökboet
      2 gold
      1 goldberg
      1 goldeagle
      2 golden
      1 golding
      1 goldmann
      1 goldstein
      1 goldtoning
      1 golf
      2 golfarmbåge
      1 golfbanor
      1 golfspelets
      1 golgi
      1 golgiapparat
      1 golgiapparaten
      1 golgiapparatens
      8 golv
      1 golvdiskmaskiner
      6 golvet
      1 golvläggare
      1 golvlister
      1 golvlyftar
      1 golvmattan
      1 golvmattor
      2 golvplattor
      1 golvvård
      1 golvvärme
      2 gom
      3 gömd
      2 gömda
      4 gömma
      1 gömmas
      4 gommen
      6 gömmer
      1 gomplastik
      2 gomseglet
      4 gomspalt
      1 gomspalter
      1 gomspenen
      1 gömställe
      2 gömställen
      1 gömt
      1 gonad
      2 gonaden
      2 gonader
      2 gonaderna
      4 gonadotropiner
      2 gonadotropinfrisättande
      1 gonadotropinnivåer
      5 gondii
      2 goniometer
      2 gonokocker
     18 gonorré
      1 gonorrheae
      1 gonorrhoea
      4 gonorrhoeae
      1 gonorrhoia
      1 gony
      1 goodman
      1 goppert
    574 gör
    285 göra
      1 göralistan
      1 göralistor
      5 göran
      1 göranden
      1 görans
     86 göras
      1 göraundvika
      1 görbersdorf
      4 gördel
      1 gördeln
      1 gördelvindlingen
      1 gördetsjälvaren
      1 gordon
      1 gore
      1 göres
      1 goretex
      1 goretexplatta
      1 gorgonen
      1 gorgoni
      1 görhåller
      1 gori
      3 gorillor
      1 görligaste
      1 göromål
    134 görs
      1 gosse
      1 gossekärlek
      3 gossen
      1 gösta
      1 göta
      1 götaland
      2 götalands
     19 göteborg
      8 göteborgs
      1 goth
      9 gotland
      1 gotlands
      1 gotländsk
      1 gotopless
      1 gotoplessorg
     45 gott
      1 gottesman
      1 gottfried
      1 gottrons
      8 gould
      1 goulds
      3 gp
      2 gproteinkopplade
      2 gps
      8 gr
     18 grå
      1 gråa
      1 graaf
      5 graafska
      3 gråaktig
      1 gråal
      1 gråblått
      1 gråbo
      2 gråbrun
      1 gråbruna
      1 gråbrunröda
    138 grad
      1 gradantal
      1 gradbeteckning
      2 grädde
      1 gräddsifoner
     31 graden
      5 gradens
     55 grader
      5 graderad
      2 graderade
      4 graderas
      1 gradering
      1 graderminut
      1 graderna
      8 graders
      1 gradienter
      1 gradindelning
      1 gradindelningen
     25 gradvis
      1 gradvisa
      2 graf
      2 grafem
      1 grafemen
      1 grafen
      3 gräfenberg
      3 grafisk
      1 grafiska
      2 grafit
      1 gråfotad
      1 grafström
      1 graftversushost
      1 grågrön
      3 grågröna
      1 grågult
      4 graham
      1 grälla
     43 gram
      1 gramfärg
      6 gramfärgning
      1 gramfärgningsresultaten
      1 graminifolius
      2 gramkg
      2 grammatik
      1 grammatiken
      1 grammatiska
      1 grammy
      4 gramnegativ
     17 gramnegativa
      1 gramnegativas
      1 grampositiv
     12 grampositiva
      1 grams
      1 gran
      1 granat
      1 granatchock
      1 granatkastare
      1 granatsplitter
      1 granbuske
      2 grand
      1 grandios
      1 grandiosa
      1 grandiositet
      1 granit
      1 graniter
      1 granlundlind
      3 grannar
      1 grannens
      2 grannländer
      9 gräns
      1 gränsar
      2 gränsdragningar
      1 gränsdragningen
     34 gränsen
      8 gränser
     10 gränserna
      1 gränsflod
      5 gränsfrekvens
      1 gränsfrekvenser
      5 granska
      5 granskade
      1 granskades
      1 granskande
      2 granskar
      3 granskas
      3 granskat
      1 granskats
      5 granskning
      1 granskningen
      1 gränslandet
      1 gränsproblematik
      1 gränssättande
      2 gränssignal
      2 gränsskikt
      1 gränsskiktet
      1 gränssnitt
      7 gränsvärde
     11 gränsvärden
      1 gränsvärdena
      6 gränsvärdet
      1 gränsyta
      1 grant
      5 granula
      1 granulär
      1 granularcellstumör
      1 granulat
      1 granulatet
      1 granulerade
      6 granulocytär
      9 granulocyter
      1 granulocytertenderar
      9 granulom
      1 granulomatos
      1 granulomatös
      1 granulomatöst
      2 granulomen
      2 granulomet
      1 granulopoes
      3 granulosaceller
      1 granulosacellerna
      1 granulosacellstumör
      1 granulosum
      2 granulosus
      1 granulum
      1 grapefrukt
      1 grapengiesser
      3 graphein
      1 grapho
      3 gråröta
      1 g�ras
      9 gräs
      1 gräsbetande
      1 gräsblad
      1 gräsgröna
      1 gräshopporna
      2 gräsmarker
      2 gräsmattor
      1 gräsrotsbyråkrat
      1 gräsrotsbyråkraterna
      1 gräsrotsrörelse
      1 grasserade
      1 grässtrån
      1 gråsvart
      3 gråt
      3 grät
      7 gråta
      1 gråtande
      1 gråtattack
      1 grateful
      4 gråter
      9 gratis
      1 gratisaffärer
      1 gratisgenerationen
      2 grått
      1 gratulationsbrev
      9 grav
     10 grava
      2 gräva
      2 gravad
      7 gravar
      1 gravare
      1 gravast
      1 grävdes
      3 gräver
      2 graves
      1 gravfältet
      1 gravfynd
     30 gravid
     56 gravida
      1 gravidaammande
      1 gravidarum
      1 gravideteter
    113 graviditet
     85 graviditeten
     12 graviditetens
     32 graviditeter
      1 graviditeterna
      1 graviditetsbevarande
     13 graviditetsdiabetes
      1 graviditetshormon
      1 graviditetshormonet
      1 graviditetshypertoni
      1 graviditetsillamående
      1 graviditetskramp
      2 graviditetslängden
      1 graviditetsmånaden
      1 graviditetsreaktion
      2 graviditetsrelaterade
      1 graviditetsstarten
      1 graviditetssymptom
      1 graviditetstalen
      3 graviditetstest
      1 graviditetstester
      1 graviditetstestet
      1 graviditetstidens
      2 graviditetstoxikos
      1 graviditetstoxikosen
      1 graviditetsultraljud
     29 graviditetsvecka
      8 graviditetsveckan
      1 graviditetsveckans
      2 graviditetsveckor
      2 graviditetsveckorna
      1 gråviolett
      1 gravis
      3 gråvit
      1 gravitationen
      1 gravkors
      2 grävling
      2 grävlingen
      2 grävlingshår
      1 grävning
      1 grävs
      1 gravsätta
      6 gravt
      1 grävt
      2 grävts
      1 gravureidoler
      7 gray
      1 grayson
      1 graziano
      2 great
      1 greater
      1 greatest
      1 greenockit
      2 greenpeace
      1 greenwalt
      1 greenwich
      1 gregorius
      1 gregory
     16 grek
      1 greken
      3 greker
      8 grekerna
      1 grekernas
      9 grekisk
    129 grekiska
      6 grekiskan
     58 grekiskans
      4 grekiske
      2 grekiskt
     23 grekland
      1 greklands
     23 gren
      1 grenad
      1 grenade
     15 grenar
      3 grenarna
      1 grenat
      4 grenen
      1 grenig
      1 greniga
      1 grenigt
      2 grenspecialitet
      2 grenspetsarna
      1 grenverket
      1 grenzschutzgruppe
      7 grepp
      2 greppa
      1 greppas
      1 greppsvaghet
      2 gres
      1 greuter
      2 grevinnan
      1 grey
      1 greyhoundhund
      1 griffeltavla
      1 grigorenko
      1 grillplatser
      1 grillspett
      3 grind
      2 grinden
      1 grinder
      1 grinig
      3 gripa
      1 gripande
      1 gripbara
      1 griper
      1 gripklor
      1 griprörelser
      1 grips
     10 gris
      8 grisar
      2 grisarna
      1 grisars
      1 grisben
      1 grisbestånd
      1 grisbetar
      1 griseus
      2 griskött
      3 grispopulationer
      1 griständer
      4 gro
      1 grobarhet
      1 grobarheten
      1 grobladsväxter
      1 gröda
      1 grodas
      1 grodben
      1 grodda
      1 groddarna
      1 groddcellstumör
      3 groddjur
      4 grodor
      7 grödor
      1 grof
      1 grogrund
      1 grohed
     16 grön
     27 gröna
      1 grönaktig
      1 grönaktiga
      2 grönalger
      1 grönblåa
      1 gröngul
      4 gröngula
      1 grönlandssäl
     23 grönsaker
      1 grönsaksblandningar
      1 grönsaksland
      1 grönsippa
      1 grönsippan
      1 grönska
      1 grönskiftande
      7 grönt
      2 grönvit
      1 grönwall
      1 groote
      3 grop
      4 gropar
      1 gropögon
      1 gror
      1 grossister
      2 grossman
      2 gröt
      2 gröten
      1 groth
      2 grotjahn
      2 grötomslag
      1 groton
      1 grötsvimmen
      1 grotta
      4 grottor
      9 group
      1 groups
      8 grov
      8 grova
      1 grovhet
      1 grovheten
      1 grovindelas
      1 grovlek
      1 grovleken
     15 grövre
      8 grovt
      1 grovtarm
      3 grovtarmen
      1 grovtarmsmynningen
      1 grovtest
      8 growth
      1 grs
      1 grubblerier
      1 grumlar
      1 grumlas
      2 grumlig
      2 grumlingar
      1 grunadare
      1 grünbaum
    536 grund
     11 grunda
      5 grundad
      9 grundade
     24 grundades
     21 grundämne
      1 grundämnen
      2 grundämnena
     10 grundämnet
      1 grundämnets
      1 grundande
      1 grundandet
      1 grundantagande
      3 grundantagandet
     14 grundar
      8 grundare
      4 grundas
      5 grundat
      1 grundats
      1 grundbehandlingen
      1 grundbetydelse
      1 grunddefinitionen
      1 grunddelar
      1 grunddemensen
      1 grundelemente
     31 grunden
      5 grunder
      1 grunderna
      1 grundexamen
      2 grundfärg
      1 grundform
      3 grundforskning
      1 grundfrekvensen
      1 grundfunktionen
      1 grundidé
      1 grundidéer
      1 grundidén
      1 grundig
      1 grundinställning
      2 grundinställningar
      2 grundkurs
      2 grundkursen
      1 grundlade
      1 grundlag
     40 grundläggande
      3 grundlig
      2 grundligt
      1 grundlinien
      1 grundlöst
      1 grundmolekyl
      3 grundnivå
      7 grundorsaken
      1 grundorsaker
      1 grundorsakerna
      2 grundprincipen
      2 grundprinciper
      1 grundrytmerna
      1 grundsärskola
      3 grundsjukdom
      1 grundskola
      2 grundskolan
      1 grundskolning
      1 grundspänning
      1 grundsteg
      1 grundstenar
      1 grundstrecken
      1 grundstreckets
      1 grundsubstans
      4 grundsubstansen
      1 grundsymptomen
      1 grundtanke
      3 grundtanken
      1 grundtillstånd
      3 grundtonen
      1 grundtoner
      1 grundtonhöjden
      1 grundtonsfrekvensen
      1 grundtyper
      4 grundutbildning
      3 grundutbildningen
      2 grundvaccination
      9 grundval
      1 grundvalen
      3 grundvatten
      1 grundversionen
      1 grünenthal
      1 grunt
    165 grupp
      1 gruppbehandling
     75 gruppen
     90 grupper
      1 gruppera
      1 grupperade
      4 grupperas
      1 grupperat
      2 grupperingar
      7 grupperna
      1 gruppers
      1 grupperspektivet
      1 gruppgäspning
      2 gruppledare
      1 gruppledarna
      1 gruppmedlemmarna
      1 gruppterapi
      1 grupptillhörighet
      1 gruppträning
      1 grupptryck
      2 grus
      1 grusade
      1 grusig
      2 gruva
      2 gruvan
      1 gruvarbetare
      1 gruvarbetet
      1 gruvdrift
      1 gruvföretagets
      1 gruvföretags
      4 gruvor
      2 grymhet
      1 grymheter
      1 grymmare
      1 grymt
      1 grymtning
      2 gryn
      1 grynig
      1 gryniga
      1 grynigheten
      1 grynigt
      1 gryta
      2 grytan
      1 grytlapp
      1 gs
      1 gsekret
      1 gsekretet
      2 gsk
      1 gsmr
      2 gte
      1 gto
      1 gtp
      1 gtphydrolys
      1 gtyp
      1 guaiacum
      1 guanin
      1 guarana
      1 guaranabär
      1 guaranin
      9 guatemala
      1 guatemalanska
      2 guayaco
      1 gubbar
      1 gubbargummor
      1 gubbegumma
     30 gud
      4 gudar
      4 gudarna
      8 guden
      2 gudinna
      2 gudinnan
      2 gudinnor
      2 gudom
      7 gudomlig
      3 gudomliga
      1 gudrun
     11 guds
      1 gudsfientliga
      2 gudstjänsten
      1 gudstjänster
      1 gudstjänstlokaler
      1 guericke
      3 guérin
      1 guidade
      3 guide
      1 guidelines
      1 guillainbarres
      2 guillainbarrés
      5 guinea
      3 guineamask
      1 guineamasken
      2 guineamaskens
      1 guineas
      4 guinness
     22 gul
     40 gula
      1 gulag
      8 gulaktig
      6 gulaktiga
      2 gulaktigt
      1 gulare
      4 gulbrun
      1 gulbruna
      1 gulbrunt
     68 guld
      2 guldaktier
      1 guldallergi
      1 gulddoublé
      1 guldgul
      1 guldgula
      1 guldhalskragar
      1 guldhalsringarna
      1 guldhalt
      1 guldkantade
      1 guldlager
      4 guldmynt
      1 guldmyntfot
      1 guldplätering
      2 guldpriset
      1 guldreserven
      2 guldskikt
      1 guldsmeder
      1 guldsmycken
      4 guldtackor
      1 guldvärdet
      1 gulesäcken
      1 gulfärga
      1 gulfärgad
      1 gulfärgat
      1 gulfärgning
      1 gulfkriget
      1 gulfkrigssyndromet
      4 gulgröna
      1 gulgrönt
      1 gulhet
      4 gulkropp
      4 gulkroppen
      1 gulkroppscysta
      1 gulkroppscystor
      3 gulkroppshormon
      1 gulkroppshormonet
      1 gullivers
      2 gullregnen
      1 gullregnsarterna
      1 gullregnsfrön
      1 gullregnssläktet
      1 gullstrand
      1 gulmarkerad
      1 guloranga
      1 gulröd
     20 gulsot
      1 gulsotsliknande
      6 gult
      1 gulvit
      3 gulvita
      2 gum
      3 gumma
      2 gummatös
      1 gummerar
     11 gummi
      1 gummiartat
      1 gummiballong
      1 gummiband
      1 gummibandsligering
      1 gummibaserade
      1 gummiboll
      1 gummicylinder
      1 gummigutta
      1 gummiinslutet
      1 gummikulor
      1 gummiliknande
      1 gummimembran
      1 gummipropp
      1 gummirankesläktet
      1 gummislang
      1 gummisula
      2 gummiträd
      2 gummor
      1 guna
      1 gunde
      1 gundishapur
      1 gundishapurakademins
      1 gungar
      1 gungflygpölar
      1 gungningar
      1 gungstolsfötter
      7 gunnar
      2 gunnarsson
      1 gunnel
      1 gunni
      1 guns
      1 gunshot
      1 guntrip
      3 gupp
      1 guppiga
      1 guppy
      1 gurgla
      1 gurgling
      1 gurion
      1 gurka
      1 gurkinläggning
      6 gurkmeja
      1 gurkmejans
      1 gurkörtens
      3 gurkväxter
      3 gustaf
      1 gustafsson
      1 gustatoriae
      5 gustav
      1 gustavsberg
      1 gustavsbergsbussen
      1 gutha
      1 guthrietest
      2 gutta
      1 guttakolhydrat
      1 guttapercha
     12 guttaperka
      1 guttaperkafallet
      1 guttaperkan
      2 guttaperkaträdet
      1 guttieballs
      3 guy
      1 guylussac
      1 guyons
      1 gvhd
      1 gwasstudie
      1 gwp
      3 gy
      1 gycklande
      1 gycklare
      1 gyges
      1 gyh
      2 gylfe
      1 gyllene
      1 gym
      1 gymnasial
      1 gymnasiala
      1 gymnasieprogram
      1 gymnasiesärskola
      1 gymnasiesärskolan
      2 gymnasieskolan
      1 gymnasieskolans
      1 gymnasiet
      1 gymnasium
      1 gymnaster
      2 gymnastik
      2 gymnastiken
      1 gymnastikövningar
      1 gymnastikskor
      1 gymnastisera
      2 gymnastiska
      1 gynecologi
      1 gynecologica
      1 gynecological
      8 gynekolog
      3 gynekologen
      5 gynekologer
      9 gynekologi
      1 gynekologiavdelningarna
      1 gynekologins
      7 gynekologisk
      1 gynekologiska
      1 gynekologmottagning
     12 gynekomasti
      4 gynna
      3 gynnar
      4 gynnas
      2 gynnat
     10 gynnsam
      8 gynnsamma
      1 gynnsammast
      8 gynnsamt
      1 gynoid
      1 győrmosonsopron
      1 gyrasproteinet
      1 gyromytrin
      1 gyron
      5 gyrus
      7 gysinge
      6 gysingevargen
      1 gysingevargens
      2 gyspergerae
      1 gyttjebaden
     50 h
    704 ha
      1 [ha]
      4 haas
      1 habenaria
      1 habenula
      2 haber
      2 haberboschmetoden
      2 habilitering
      1 habiliteringsenhet
      1 habiliteringshund
      1 habiliteringshundar
      2 habiliteringshunden
      1 habiliteringshundens
      1 habiliteringshundlegitimationen
      1 habiliteringshundutbildning
      3 habit
     11 habitat
      1 habitatet
      1 habitatförlust
      1 habituell
      1 habitueras
      2 habituering
      3 haccp
      2 hace
      1 häckar
      1 hacken
      1 hackigt
      1 hackor
      1 häda
      2 hädanefter
    434 hade
      1 hades
      1 hädiskt
      1 hadrianus
      1 haematologisten
      1 haematomyzus
     10 haemophilus
      1 haemosideros
    115 haft
      1 häftämne
      2 häftig
      3 häftiga
      5 häftigt
      1 häftplåster
      1 hagalund
      3 hagalunds
      2 hagar
      1 hagen
      1 håglös
      1 hagtorn
      8 hahnemann
      3 hahnemanns
      1 haida
      1 haima
      1 haimorrhois
      3 haiti
      1 haja
      1 hajar
      1 hajen
      2 hajj
      1 hajk
      5 haka
      2 hakade
      5 hakan
      2 håkansson
      4 hakar
      1 hakarna
      1 hakat
      1 hakmask
      1 häkta
      1 hal
     33 hål
      1 häl
      2 hala
      2 håla
      1 halabja
      1 halal
      1 hälar
      3 hälbenet
      1 haldane
      2 haldaneeffekten
      3 haldol
      1 haldolbehandling
      1 haldols
      1 hålen
      8 hälen
      8 hålet
      1 halford
      1 hålförstärkning
      1 hålfot
      1 hålfotsinlägg
      6 hälft
     88 hälften
      1 halglatt
      1 halidjoner
      4 hålighet
      1 håligheten
      6 håligheter
      1 håligheterna
      1 haliotissnäckan
      1 halit
      1 halka
      1 halkade
      1 hall
     55 håll
    125 hålla
      4 hälla
      5 halland
      1 hållande
      2 hallands
      2 hallandsåsen
      3 hållare
     17 hållas
      2 hällas
      4 hållbar
      1 hällbär
      3 hållbara
      2 hållbarhet
      3 hållbarheten
      1 hållbarhetsskäl
      1 hållbarhetstid
      3 hållbarhetstiden
      2 hållbart
      1 hällde
      1 hälldes
      1 halleffekten
      1 hållen
     82 håller
      1 häller
      1 hallersteinii
      1 hålles
     15 hållet
      1 hållfasthet
      6 hållit
      2 hållits
      3 hållna
     12 hållning
      2 hållningen
      1 halloffamebasebollspelaren
      2 hallon
      2 hällristningar
     32 hålls
      1 hällts
     11 hallucination
      1 hallucinationen
     72 hallucinationer
     11 hallucinationerna
      1 hallucinatus
      1 hallucinera
      2 hallucinerar
     12 hallucinogena
      8 hallucinogener
      1 hallucinogent
      2 hallucinoser
      2 haloalkan
      1 haloalkaner
      1 haloform
      3 halogenalkan
      1 halogenatom
      1 halogener
      2 halogenerad
      1 halogenerade
      1 halogenering
      1 halogeniseras
      1 halogenlampa
      1 halogenlampor
      1 halogentyp
      4 hålor
      8 halotan
      1 halothan
      3 hålrot
     12 hålrum
      1 hålrummen
      3 hålrummet
      1 hålrummets
      1 hålrumssystem
     11 hals
    154 hälsa
      1 hälsades
     33 hälsan
      2 hälsans
      1 hälsaohälsa
      1 halsartärer
      1 halsartärerna
      3 halsband
      4 halsbränna
      1 halsbrännaoch
      1 halsdoktor
      1 halsduk
      1 halsdukar
     48 halsen
      1 hälsena
      1 hälsenan
      1 hälsenesnitt
      5 halsens
     15 halsfluss
      1 halsgropen
      2 halshuggning
      2 halsinfektion
      1 halsinfektioner
      1 halsinflammation
      1 hälsingland
      1 hälskål
      1 halskota
      1 halskotpelaren
      1 halslymfknutor
      1 halsmandelsstenar
      2 halsmandelvecken
      1 halsmandlar
      7 halsmandlarna
      4 halsmandlarnas
      1 halsmuskulaturen
      2 hälsning
     47 hälso
      2 hälsoaspekter
      5 hälsobefrämjande
      2 hälsobegrepp
      2 hälsobegreppet
      3 hälsobokslut
      2 hälsobokslutet
      4 hälsobringande
      2 hälsocentral
      1 hälsodataregister
      1 hälsodebatten
      3 hälsodefinition
      1 hälsodefinitionen
      1 hälsodefinitioner
      1 hälsodeklaration
      2 hälsodepartement
      1 hälsodryck
      1 hälsoeffekt
     16 hälsoeffekter
      2 hälsoekonomi
      2 hälsoekonomiska
      1 hälsoenkät
      1 hälsoentrepenören
      5 hälsofara
      1 hälsofaran
      3 hälsofarliga
      2 hälsofaror
      2 hälsofarorna
      1 hälsofördelar
      6 hälsofrämjande
      1 hälsogrundade
      1 hälsoit
      1 hälsojournalisten
      2 hälsokonsekvenser
      1 hälsokontorets
      1 hälsokontroll
      3 hälsokontroller
      1 hälsokontrollerna
      2 hälsokost
      2 hälsokostaffärer
      1 hälsokostbutiker
      1 hälsokostsammanhang
      1 hälsolevernet
      1 hålsöm
      1 hälsomässig
      1 hälsomässiga
      1 hälsomat
      1 hälsominister
      2 hälsoministeriet
      2 hälsoministrar
      1 halsområdet
      1 hälsomyndighet
      1 hälsomyndigheter
     13 halsont
      6 hälsooch
      1 hälsopåverkan
      2 hälsoperspektiv
     18 hälsoproblem
      1 hälsoprodukt
      6 hälsoprogram
      1 hälsoprogrammen
      1 hälsorelaterad
      1 hälsorelaterade
      1 hälsoriktig
      7 hälsorisk
     18 hälsorisker
      2 hälsoriskerna
      9 hälsosam
      5 hälsosamma
      1 hälsosammare
      9 hälsosamt
      2 hälsoskadliga
      7 hälsoskäl
      1 hälsoskydd
      1 hälsosvikt
      9 hälsotillstånd
      3 hälsotillståndet
      1 hälsoupplysning
      4 hälsovådliga
      2 hälsovådligt
      7 hälsovård
      1 hälsovårdande
      3 hälsovården
      1 hälsovårdsarbete
      1 hälsovårdsdepartementet
      1 hälsovårdslära
      1 hälsovårdsministreriet
      1 hälsovårdsmyndigheterna
      1 hälsovårdspersonal
      7 hälsporre
      2 hälsporren
      1 halspulsådern
      2 halsregionen
      1 halsring
      5 halsringar
      1 halsryggen
      1 halssjukdomar
      1 halsskrofler
      1 halsspecialisten
      1 halstablett
      8 halstabletter
      1 halsvenstas
     24 halt
      1 halta
      3 hälta
      2 håltagning
      1 håltagningar
      1 håltagningen
      1 haltande
     24 halten
     46 halter
      8 halterna
     12 halv
     11 halva
      1 halvädelstenar
     14 halvan
      1 halvannat
      3 halvår
      2 halvåret
      3 halvårs
      1 halvårslinser
      1 halvårsvis
      2 halvautomatiska
      1 halvbad
      2 halvbror
      1 halvbrors
      1 halvcirkel
      1 halvcirkelformad
      1 halvcirkelns
      5 hålvenen
      1 hålvener
      1 hålvenerna
      2 halvera
      1 halverades
      2 halveras
      2 halverats
      9 halveringstid
      4 halveringstiden
      1 halveringstider
      1 halvfasta
      2 halvfullt
      1 halvgudomlig
      1 halvkloten
      6 halvklotet
      1 halvklotets
      1 halvklotformigt
      1 halvknuten
      1 halvkupor
      1 halvlåg
      1 halvledare
      1 halvligga
      1 halvliter
      1 halvmåne
      1 halvmåneformad
      1 halvmåneformig
      1 halvmetall
      1 halvmetalliskt
      2 halvön
      1 halvöppna
      1 halvor
      1 halvorna
      2 halvsides
      1 halvsidig
      1 halvsidiga
      1 halvsittande
      1 halvskugga
      1 halvskuggig
      1 halvslutna
      1 halvsovande
      1 halvstrukturerade
      1 halvsyntetiskt
      5 halvt
      1 halvterminskurser
      1 halvtidspausens
      1 halvtidsuppträdandet
      1 halvtimma
      7 halvtimme
      2 halvtomt
      1 halvtorra
      1 halvvägsboende
      1 ham
      1 hamam
      4 hamartom
      1 hamartomet
      1 hamilton
      1 hamlet
     23 hämma
      4 hämmad
      5 hämmade
     10 hämmande
     45 hämmar
      1 hammarberg
      2 hammare
      1 hämmare
      1 hammaren
      7 hämmas
      5 hämmat
      1 hammer
      4 hamn
     11 hamna
      2 hamnade
     34 hamnar
      1 hämnas
      6 hamnat
      3 hämnd
      1 hämndmotiv
      2 hamnen
     11 hämning
      1 hämningar
      1 hämningen
      1 hämningsdepressioner
      1 hämoglobin
      1 hampa
      1 hampafrön
      1 hams
      1 hamster
      2 hamstrar
      1 hamsun
      3 hämta
      6 hämtad
      6 hämtade
      3 hämtar
      6 hämtas
      4 hämtat
      2 hämtats
      1 hämtplats
      1 hamul
    449 han
      2 hån
      7 hanar
      1 hånar
      6 hanarna
      3 hanblommor
      2 hanblommorna
    144 hand
     15 hända
      1 handaggregat
      2 handakupunktur
      1 handalfabet
      1 handanlag
      1 hand�armvibrationssyndrom
      2 handboken
      1 handdarrningar
      1 handdesinfektion
      1 handdesinfektionsmedel
      2 handdisk
      1 handdiskas
      1 handdrivna
      8 handduk
      7 handdukar
      4 handduken
      1 handdukens
      1 handduksdagen
      1 handdukstorkar
      1 handdukstorkas
      1 handduksväv
      1 handduschar
      4 hände
      1 handeksem
     10 handel
     11 handeln
      1 handelsbalansen
     12 händelse
      4 händelseförlopp
      2 händelseförloppet
      1 händelsekedja
      1 händelsekedjan
     11 händelsen
     33 händelser
      4 händelserna
      1 händelserssjukdomarsföreteelsers
      1 handelsfartyg
      1 handelsgödsel
      1 handelsknutpunkt
      1 handelsknutpunkterna
      3 handelsmän
      6 handelsnamn
      2 handelsnamnen
      4 handelsnamnet
      1 handelspolitik
      2 handelspost
      1 handelsstaden
      1 handelstillgängligt
      2 handelsvägar
      1 handelsvara
      1 handelsvaran
      1 handelsvaror
      1 handelsvillkor
     34 handen
      7 handens
     73 händer
      1 händerarmar
      1 händerfingrar
     45 händerna
      1 händernas
      1 händervid
      1 handfängsel
      2 handfat
      2 handflata
      5 handflatan
      4 handflator
      5 handflatorna
      3 handflikiga
      1 handfull
      1 handgranat
      2 handgrepp
      1 handgreppet
      1 handgripliga
      2 handhaft
      3 handhar
      1 handhas
      3 handhavande
      5 handhygien
      1 handicare
      1 händighetsstörningar
     24 handikapp
      1 handikappad
      1 handikappade
      5 handikappande
      1 handikappbegreppet
      1 handikappet
      1 handikappförbunden
      1 handikappförening
      1 handikapporganisation
      1 handikapporganisationer
      1 handikapptoaletter
      2 handikappvetenskap
      1 handjur
      1 handkirurg
      2 handkirurgi
      1 handkontrollen
      1 handkontroller
      1 handkontrollerna
      2 handkraft
      1 handkrämer
     25 handla
      6 handlade
      1 handläggaren
      1 handlägger
      3 handläggning
      1 handläggningen
      1 handläggs
      8 handlande
     91 handlar
      1 handlas
      4 handlat
      2 handled
      4 handleda
      3 handledare
      1 handledaren
      1 handledd
     11 handleden
      1 handledens
      3 handleder
      1 handlederna
      4 handledning
      1 handledsortoser
      1 handledsskärandesyndrom
      1 handledsskena
      1 handlexikon
      1 handlin
     14 handling
     39 handlingar
     13 handlingen
      1 handlingsförlamning
      4 handlingsförmåga
      1 handlingsinriktning
      1 handlingslinje
      1 handlingsmönster
      1 handlingsplan
      3 handlingsplanen
      1 handlingsplaner
      1 handlingsprogrammet
      1 handlingsrelaterad
      1 handlingssättet
      2 handlingsutrymme
      1 handmotorikcentra
      6 handpåläggning
      1 handrörelser
      2 handrullade
      1 handrullning
      4 hands
      1 handsaker
      2 handskar
      5 handskas
      1 handsken
      1 handskrifter
      1 handslag
      9 handsprit
      1 handspriten
      1 handsprithanddesinfektion
      1 handstycket
      9 handtag
      1 handtagen
      5 handtaget
      1 handtagets
      2 handtork
      1 handtremor
      7 handtvagning
     12 handtvätt
      2 handtvättningen
      6 hane
     10 hanen
      2 hanens
      1 hanfisk
      1 hänföra
      5 hänföras
      1 hänförd
      3 hänförs
     12 hänga
      2 hangametofyten
      6 hängande
      2 hängas
      4 hängde
     31 hänger
      1 hängfuchsia
      1 hängighet
      1 hängigt
      2 hängiven
      1 hängivenhet
      1 hängivet
      1 hängivit
      1 hänglobelia
      3 hängning
      2 hängs
      2 hängt
      2 hängtorka
     13 hanhon
      1 hanindivider
      1 hankön
      1 hankottarna
      2 hanlarver
      1 hanlig
      5 hanliga
      1 hanligt
      1 hanmaskar
      3 hann
      1 hannah
      7 hannar
      5 hannarna
      1 hannarnas
      2 hanne
      4 hannen
      1 hannens
      1 hannibal
      1 hanÖ
      2 hanorganet
      1 hanplantan
      1 hanplantor
    130 hans
      1 hansans
      5 hänseende
      1 hänseenden
      2 hansen
      4 hansens
      1 hansheinrich
      2 hanshennes
      1 hansletsgräs
      1 hansson
      1 hansurta
      1 hänsyftning
     32 hänsyn
      1 hänsynslösa
      1 hänsynslöshet
      5 hänt
      1 hantaanvirus
      1 hantan
      3 hantavirus
     72 hantera
      2 hanterades
      1 hanterande
     14 hanterar
     20 hanteras
      2 hanterat
      1 hanterats
      1 hanterbar
      1 hanterbara
      7 hanterbarhet
      1 hanterbart
     16 hantering
      7 hanteringen
      1 hanterlig
      1 hanterliga
      1 hanterligt
      3 hantverkare
      1 hantverkartradition
      1 hantverksmässiga
      2 hantverksmässigt
      1 hantverksorganiserade
      1 hanvaran
      2 hänvisa
      2 hänvisade
     11 hänvisar
      2 hänvisas
      1 hänvisat
      6 hänvisning
      1 haparanda
      4 hape
      3 haploid
     11 haploida
      1 haplotypen
      1 häpnadsväckande
      2 hapten
      4 haptoglobin
      1 hapy
   5291 har
     56 hår
    183 här
      1 häradet
      1 häradsrätten
      2 harald
      5 harar
      1 hararna
     18 håravfall
      2 håravfallet
      1 hårbärande
      1 härbärgen
      1 härbärgera
      1 harbeståndet
      1 harbor
     11 hårborttagning
      1 hårborttagningskräm
      1 hårborttagningsmetod
      8 hårbotten
      1 hårbottnen
      1 harbour
      3 hårceller
      5 hårcellerna
      1 hårcellsleukemi
     38 hård
     20 hårda
      2 härdar
     12 hårdare
      1 härdas
      1 hårdast
      2 härdat
      1 hårdbevakad
      1 härden
      1 hårdgummi
      1 hårdheten
      2 härdig
      1 härdiga
      1 härdighet
      1 hardjur
      1 hårdkokta
      1 hårdnad
      2 hårdnar
      2 hardness
      1 härdning
      1 härdningsprocess
      1 härdningsprocessen
      3 hårdost
      1 hårdostar
      1 hårdplast
      1 härdplast
      1 härdplaster
      1 hårdrocksbandet
      1 hårdröntgenstrålning
      1 hårdträna
      3 hårdvara
      1 hårdvävnad
      4 hare
      3 harem
      1 haremsdamer
      5 håren
      3 hares
     27 håret
      1 hårfagers
      2 hårfärg
      3 hårfärger
      1 hårfärgningsmedel
      1 hårfärgsprodukter
      1 hårfästet
      1 hårfolliklar
      1 hårfön
      1 härförs
      1 hårgurkssläktet
      1 häri
      4 härifrån
     12 hårig
      4 håriga
      1 hårigt
      6 härjade
      2 härjar
      2 härjat
      2 härjningar
      1 harkla
      2 harklar
      1 harklingar
      1 hårklippning
      3 härkomst
      1 härkomster
      1 hårkors
      1 hårkvalitet
      4 härleda
     10 härledas
      1 härleder
      1 härledning
      1 härledningen
      3 härleds
      2 härlett
      1 hårliknande
      1 hårlösa
      1 hårlyft
      3 harm
      4 härma
      1 harman
      2 härmar
      3 härmed
      1 hårmedel
      3 harmlösa
      3 harmlöst
      1 härmningar
      3 harmoni
      1 harmonisk
      2 harmoniska
      1 hårnålar
      1 härochnuvarande
      1 harold
      6 harpest
      1 hårpreparat
      1 harpuner
      1 hårredskap
      1 hårreducering
      1 harrelson
      1 hårremmen
      1 harriet
      2 harrison
      1 hårrör
     19 härrör
      1 härröra
      2 härrörande
      1 härrörde
      1 hårrötter
      3 harry
      2 hårsäck
      8 hårsäckar
      5 hårsäckarna
      2 hårsäckarnas
      3 hårsäcken
      4 hårsäcksgrupper
      1 hårsäcksinflammation
      2 hårsäcksinflammationer
      1 hårsäckssjukdom
      1 hårsäckstransplantat
      3 härskare
      1 härskat
      1 härskna
      1 härsknar
      1 härskning
      2 härstamma
      1 härstammade
      1 härstammande
     34 härstammar
      1 härstamning
      4 hårstrå
      6 hårstrået
      9 hårstrån
      6 hårstråna
      1 hårstrår
     56 hårt
      1 härtåg
      1 hartdegen
      4 hartelius
      1 harter
      3 hartmann
      3 hårtransplantation
      1 hårtransplantationsmetoder
      2 harts
      4 hartser
      1 hartset
      1 hartskloroform
      2 hårtvätt
      1 hårtvättar
      1 hårtvätten
      1 hårtyper
      1 härutöver
      1 härva
      1 hårvårdsprodukt
      2 hårvårdsprodukter
     10 hårväxt
      5 harvey
      7 härvid
      2 has
      1 hasande
      7 hasardspel
      2 hasardspelsyndrom
      3 hashimotos
      1 hassan
      1 hasselakollektivet
      1 hasselbalch
      2 hasselnötter
      1 hasselnötterparanötter
      1 hasselström
      1 hasslerianus
     10 häst
     39 hästar
      1 hästarbr
      1 hästarna
      1 hästbane
      1 hästdjur
      1 hästen
      1 hästfibbla
      2 hästfluga
      1 hästflugan
      1 hästhår
      3 hästhov
      1 hästhovar
      1 hästhovens
      1 hästhovsört
      5 hastig
      3 hastiga
     28 hastighet
      6 hastigheten
      4 hastigheter
      1 hastighetsbegränsning
      1 hastighetsbestämmande
      1 hastighetsgränsen
      1 hastighetsuppgifterna
     19 hastigt
      1 hastings
      1 hästkadaver
      1 hästkastanj
      2 hästmedicin
      1 hästsjukdomar
      1 hästsko
      2 hästskoformade
      2 hästskonjure
      1 hästskötsel
      2 hat
      3 hata
      1 hatbrott
      1 hatha
      8 hathayoga
      1 hatschek
      1 hätsk
      7 hatt
      1 hätta
      1 hattar
      1 hattdiameter
      6 hatten
      2 hattens
      1 hatter
      1 hattformen
      1 hatthuden
      3 hattmakare
      1 hatton
      1 hattsvamparna
      1 haung
      1 haurio
      1 hauser
      1 haustor
      1 haustorialhyfer
      3 haustorier
      1 haustorierna
      1 haustra
      1 haustrierna
      1 haute
      1 haüy
      6 hav
      4 häva
      3 havande
      2 havandeskap
      2 havandeskapet
      2 havandeskapsdiabetes
      6 havandeskapsförgiftning
      1 hävas
      2 hävd
      6 hävda
     12 hävdade
     47 hävdar
      3 hävdas
      6 hävdat
      2 hävdats
      1 have
      1 häver
      1 havererar
      1 haveriet
     16 havet
      1 havorringen
      5 havre
      1 havregryn
      1 havregurtsoygurt
      1 havremjölk
      3 havrix
      2 havs
      3 hävs
      1 havsbotten
      1 havsbottnen
      3 havsgeting
      4 havsgetingen
      1 havsgetingens
      1 havsnära
      1 havsnivå
      2 havsormar
      1 havsormarna
      1 havsörnen
      3 havssalt
      3 havsskada
      1 havssköldpaddor
      1 havsskummet
      1 havsstränder
      1 havstränder
      1 havstulpaner
      1 havsvågor
      7 havsvatten
      1 havsvattennivån
      1 havsvindar
      1 hawaii
      1 hawaiiansk
      1 hawaiianskt
      1 hawkins
      4 häxeri
      3 häxkonsten
      1 häxkonstnärer
      3 häxkvast
      1 häxmästare
      1 häxmjölk
      6 häxor
      6 häxorna
      1 häxornas
      1 häxringar
      2 häxsabbat
      2 häxsabbater
      1 häxsalva
      1 häxsalvor
      1 hazard
      2 hazell
      3 hb
      1 hblockerare
      1 hbo
      1 hbobehandling
      1 hbon
      7 hbov
      1 hbtnormen
      1 hbvärde
      1 hc
      3 hcc
      4 hcg
      1 hcgnivån
      6 hcl
      2 hco
      1 hcov
      1 hcp
      2 hcrtorexin
      2 hd
      1 hdl
      1 hdlkolesterol
      1 hdp
      1 headache
      2 headings
      2 healern
     10 healing
      1 healingbehandling
      1 healingen
      1 healningar
     31 health
      2 healthcare
      1 hearing
      5 heart
      1 heartbrand
      1 heartbrandmärkningen
      1 heat
      1 heatrepetitioner
      3 heavy
      1 hebamme
      1 hebe
      3 hebefren
      1 hebosteotomi
      1 hebreiska
      1 hedar
      1 hedén
      1 heder
      1 hederacae
      1 hedern
      1 hederskors
      2 hederstitel
      2 hedge
      1 hednisk
      2 hedoni
      1 hedonistisk
      2 hedra
      2 hedrar
      1 hegel
      1 heidenstam
      1 heimlich
      1 heimlichmanövern
      3 heinrich
      1 heinz
      1 heittää
      2 hej
      5 hejda
      1 hejdade
      2 hejdar
      2 hejdas
      1 hektakomber
      2 hektar
      1 hekton
     33 hel
    342 hela
      1 helades
      1 helägt
     10 helande
      1 helandets
      1 helar
      1 helautomatiska
      2 helblod
      1 helbräddade
      1 helbrägda
      1 helcellsvaccin
      1 helen
      1 helena
      1 helgat
      1 helgeandshus
      1 helgedomar
      2 helgon
      1 helgonet
      1 helgonkult
     14 helhet
      1 helheten
      2 helhetsförståelse
      1 helhetsperspektiv
      1 helhetssyn
      1 helichrysum
      5 helicobacter
      3 helig
      7 heliga
      7 helige
      1 heliges
      1 helighet
      1 heligt
      1 helikal
      1 helikopterexpedition
      2 helikoptrar
      2 helios
      1 heliox
      4 helium
      2 helix
      1 �helixdomäner
      1 helixen
      1 helkonstigt
      1 helkroppsdatortomografi
      1 helkroppspletysmograf
      1 helkroppsreflexen
      1 helkroppsröntgen
      1 helkroppsvibrationer
      1 hell
      2 helleborus
      1 helleboruskur
      1 hellenistiska
     94 heller
      1 hellered
      1 hellers
      1 hellmut
      1 hellmuth
      1 helloweenbrian
      1 hellp
      4 hellre
      1 helmholtz
      1 helmut
      5 heloderma
      2 helosan
      1 helping
      1 helsilikonkateter
      1 helsilikonkatetrar
      2 helsingborg
      7 helsingfors
      1 helsingforsdeklarationen
     64 helst
      1 helsvart
      1 helsydda
      1 helsyskon
    336 helt
      4 heltäckande
      1 heltid
      1 heltidsanställd
      3 heltidsstudier
      1 heltidstjänster
      1 helvegetarisk
      2 helveteseld
      3 helvetet
      2 helvit
      2 helvita
     54 hem
      3 hemagglutinin
      1 hemangiom
     18 hemangiosarkom
      1 hemangiosarkomet
      1 hemanvändare
      1 hematemes
      1 hematochezi
      1 hematokezi
      2 hematokrit
      3 hematologi
      2 hematologin
      1 hematologins
      1 hematologiska
      1 hematom
      1 hematopoes
      2 hematopoesen
      1 hematopoetisk
      2 hematopoetiska
      1 hematospermi
      6 hematuri
      1 hematurikateter
      1 hematurikatetrar
      5 hembehandling
      1 hembehandlingpatienten
      6 hembesök
      1 hemdammsugare
      1 hemdelar
      1 hemelektronik
      1 hemfärden
      1 hemfödd
      1 hemfödslar
      1 hemföll
      3 hemförlossning
      3 hemförlossningar
      1 hemgång
      1 hemgjorda
      4 hemgrupp
      3 hemgruppen
      1 hemgruppens
      2 hemianopsi
      1 hemingway
      1 hemingways
      2 hemipares
      1 hemipenisar
      4 hemipterus
      2 hemisfär
      5 hemisfären
      4 hemisfärotomi
      2 hemjärnet
      1 hemklinik
      1 hemkommande
      1 hemkommen
      1 hemkomst
      2 hemland
      2 hemlandet
      2 hemläxor
      1 hemlichmanövern
      2 hemlig
      3 hemliga
      3 hemlighet
      1 hemligheten
      1 hemligheter
      1 hemlighetsmakeriet
      2 hemligt
      1 hemlinjen
      1 hemlösa
      1 hemlöshet
     27 hemma
      7 hemmabruk
      1 hemmadialyserande
      2 hemmafixare
      3 hemmagjord
      1 hemmagjorda
      1 hemmahamnen
      1 hemmahörande
      1 hemmamamma
      2 hemmasittare
      1 hemmawarande
      2 hemmen
     23 hemmet
      1 hemmetpå
      1 hemmets
      2 hemmiljö
      1 hemmiljön
      1 hemmorragisk
      1 hemoblogin
     14 hemodialys
     16 hemofili
      1 hemofobi
     45 hemoglobin
      1 hemoglobiner
     18 hemoglobinet
      9 hemoglobinets
      1 hemoglobinkomplexet
      2 hemoglobinkoncentrationen
      2 hemoglobinmolekyl
      4 hemoglobinmolekylen
      1 hemoglobinmolekylerna
      1 hemoglobinsjukdomar
      1 hemoglobinsyntes
      2 hemoglobinsyntesen
      1 hemokoncentration
      4 hemokromatos
      8 hemolys
      1 hemolyserar
      1 hemolysis
      3 hemolytisk
      2 hemolytiska
      4 hemoptys
      1 hemorragi
     15 hemorragisk
      1 hemorrhagic
      1 hemorrhoid
      3 hemorrojd
      2 hemorrojdala
      1 hemorrojdektotomi
     35 hemorrojder
      2 hemorrojderna
      2 hemorrojdoperation
      3 hemorrojdplexus
      1 hemorrojdsmärta
      1 hemorrojdsymtom
      2 hemort
      4 hemostas
      5 hemostasen
      1 hemostasens
      2 hemotoxin
      1 hemotoxiner
      1 hemprotein
      1 hemresan
      3 hemsida
      1 hemsjukvård
      2 hemsjukvården
      1 hemska
      1 hemskheter
      1 hemskt
      1 hemsökte
      1 hemsöktes
      1 hemtextilier
      2 hemtjänst
      7 hemtjänsten
      1 hemtjänstgrupp
      1 hemtjänstpersonalen
      4 hemtjänstutförare
      1 hemuppgift
      1 hemvård
      2 hemvården
      1 hemvårdens
      1 hemvist
      1 hemwist
      1 hen
      1 henbane
      2 henderson
      1 hendersonhasselbalchekvationen
      1 hendrix
      3 henna
     15 henne
     44 hennes
      1 henning
      1 henosis
      3 henri
      1 henrialexandre
      1 henrietta
      4 henrik
      6 henry
      2 hensbroek
      1 henschen
      1 hep
      2 hepafilter
      5 heparin
      1 heparinbehandling
      2 hepatica
      3 hepaticus
      1 hepatikus
      2 hepatis
      1 hepatisk
      1 hepatiskt
     79 hepatit
      1 hepatitis
      1 hepatitsmitta
      1 hepatitsymptom
      1 hepatitvirus
      2 hepatocellulär
      1 hepatocellulärt
      2 hepatocyter
      4 hepatocyterna
      1 hepatologin
      1 hepatom
      2 hepatomegali
      1 hepatopancreaticasphincter
      5 hepatosplenomegali
      1 hepatotoxin
      1 hepburn
      1 heppenheim
      3 heracleum
      1 heraldiken
      1 heraldiskt
      2 herba
      6 herbert
      1 herbicid
      2 herbicider
      1 herbivorer
      1 herdecke
      1 herdefolk
      1 hereditär
      3 hereditärt
      2 hereditet
      1 heringbreuereffekten
      1 heringbreuerreflexen
      1 heringbreuers
      1 hermafrodism
      1 hermafrodit
      2 hermafrodita
      3 hermafroditer
      2 hermafroditiska
      3 herman
      1 hermandad
      5 hermann
      1 hermelin
      1 herminie
      1 hernia
      1 hernierar
      1 herniering
      2 hero
      2 herodotos
      1 heroic
      5 heroin
      1 heroiska
     12 herpes
      1 hérpes
      1 herpesblåsor
      1 herpessjukdom
      5 herpesvirus
      1 herpositivitet
      2 herptiler
      1 herr
      2 herrar
      1 herrbågar
      1 herrefolk
      1 herrens
      4 herrgård
      2 herrnstein
      1 herrparfym
      3 hertz
      1 hervey
      2 herxheimers
      4 hes
      1 heselden
      8 heshet
      1 hesheten
      1 hesketh
      2 hesron
      1 hesyre
      6 het
      4 heta
     50 heter
      2 hetero
      1 heteroanamnes
      1 heterocyklisk
      1 heterocykliska
      1 heterogen
      1 heterogenitet
      1 heterogent
      6 heterokromi
      7 heterosexuella
      2 heterosexuellt
      1 heterotropiskt
      3 heterozygot
      1 heterozygota
      2 hetsat
      1 hetsätning
      1 hetsen
      1 hetsiga
      5 hett
      8 hetta
      1 hettade
      3 hettan
      2 hettar
      3 hettas
      6 hette
      1 heu
      1 heverteffekten
      1 hewson
      1 hexabutyldistannan
      1 hexameter
      1 hexametylentetramin
      1 hexeditin
      1 hexenuronsyra
      1 hexis
      1 hexogen
      1 hf
      3 hfa
      3 hg
      1 hgjoner
      1 hgs
      3 hhs
      1 hi
      1 hiaa
      2 hiatusbråck
      1 hibernal
      1 hibernalet
      1 hibvaccinet
      1 hielpa
      1 hiemalis
      1 hiemis
      1 hierarki
      1 hierarkin
      1 hierarkisk
      1 hierarkiska
      1 hierosolymitanus
      6 high
      1 highaltitude
      3 highly
      2 highway
      1 higoumenakis
      1 hijras
      5 hikikomori
      1 hikikomorí
      4 hikikomorier
      4 hikikomorierna
      1 hikikomoriernas
      2 hildebrand
      1 hildegard
      2 hill
      1 hillman
      1 hiltons
      1 hiltula
      2 himalaya
      5 himlen
      1 himmel
      2 himmelen
      1 himmelriket
      1 himmelsk
      1 himmerfjärdsverket
      1 himmler
     14 hinder
      1 hinderbana
      1 hindi
      1 hindins
     41 hindra
      2 hindrade
      1 hindrades
      1 hindrande
     42 hindrar
      9 hindras
      1 hindrat
      5 hindret
      1 hindu
      3 hinduer
      1 hinduisk
      2 hinduiska
      2 hinduism
     10 hinduismen
      3 hinduismens
      1 hinduistiska
      6 hindustan
      1 hingstar
      2 hink
     13 hinna
      1 hinnan
     21 hinner
      1 hinnliks
      2 hinnor
      1 hinnorna
      1 hinz
      1 hinzii
      1 hippie
      2 hippies
      1 hippobosca
      2 hippoboscidae
     27 hippocampus
      1 hippocampusstrukturen
      2 hippocrates
      3 hippocraticum
     18 hippokrates
      2 hippokratiska
      1 hiprex
      1 hiragana
      2 hirs
      4 hirsutism
      1 hirticarpus
      1 hirudin
      2 hirudo
      1 his
      2 hisa
      3 hiss
     25 histamin
      1 histamine
      1 histaminer
      2 histidin
      1 histidingruppernas
      1 histidinresternas
      1 histocompatibility
      1 histokompatibilitetsantigen
      1 histokompatibilitetskomplex
      2 histologi
      1 histologin
      3 histologisk
      4 histologiska
      2 histologiskt
      1 histoner
      2 histoplasma
      2 histoplasmos
    156 historia
     15 historien
      6 historiens
      6 historier
      2 historierna
      2 historieskrivning
     64 historik
      3 historiken
      1 historikern
      7 historisk
     19 historiska
     32 historiskt
      2 history
      2 histrionisk
     11 hit
      1 hitchcock
      1 hitchcockianus
      1 hitintills
      3 hitler
      1 hitlers
     74 hitta
     11 hittade
     13 hittades
     18 hittar
     25 hittas
     16 hittat
     11 hittats
     15 hittills
     83 hiv
     12 hivaids
      1 hivassocierad
      1 hivassocierade
      1 hivb
      1 hivbehandling
      1 hivbromsmediciner
      1 hivepidemins
      1 hivförekomsten
      1 hivinfekterad
      2 hivinfekterade
     12 hivinfektion
      2 hivinfektionen
      1 hivnegativa
      4 hivöverföring
      4 hivpositiv
     10 hivpositiva
      1 hivrelaterade
      1 hivsmitta
      6 hivsmittade
      1 hivsmittan
      1 hivsmittat
      1 hivstammar
      1 hivtesten
      2 hivvirus
      4 hivviruset
      2 hjälm
      2 hjalmar
      3 hjälmar
      1 hjälmars
      1 hjälmbönssläktet
      2 hjälmen
      1 hjälmformigt
      1 hjälmmössa
    376 hjälp
     64 hjälpa
      1 hjälpämnen
      1 hjälpämnet
      2 hjälpande
      1 hjälpare
      1 hjälpas
      1 hjälpbehovet
     12 hjälpen
      1 hjälpenbehandling
      1 hjälpenlådor
     76 hjälper
      1 hjälpligt
      1 hjälplösa
      1 hjälplöshet
     66 hjälpmedel
      1 hjälpmedelscentral
      1 hjälpmedelsindustri
      1 hjälpmedelsinstitutet
      2 hjälpmedlen
      1 hjälporganisationer
      1 hjälps
      1 hjälpsamt
      7 hjälpt
      4 hjälpta
      7 hjälpte
      1 hjälpverktyg
      1 hjältar
      1 hjältarnas
      3 hjälte
      1 hjältefigur
      1 hjältemodiga
      2 hjältinnor
      2 hjälv
      1 hjärn
     25 hjärna
      1 hjärnaktivering
      2 hjärnaktivitet
      1 hjärnaktivitetsnivåer
    307 hjärnan
     65 hjärnans
      1 hjärnartären
      1 hjärnavbildningstekniker
      1 hjärnbark
     20 hjärnbarken
      2 hjärnbarkens
      1 hjärnbarksneuron
     16 hjärnblödning
      1 hjärnblödningar
      1 hjärnblödningarna
      6 hjärnbryggan
      5 hjärnceller
      1 hjärncellerna
      2 hjärncentra
     10 hjärndöd
      1 hjärndöda
      1 hjärndödsdiagnostik
      1 hjärnfel
      1 hjärnförändringar
      1 hjärnfunktion
      2 hjärnfunktioner
      1 hjärnfunktionerna
      5 hjärnhalva
      5 hjärnhalvan
      1 hjärnhalvorna
      1 hjärnhandikapp
      2 hjärnhinna
      7 hjärnhinnan
      4 hjärnhinne
     23 hjärnhinneinflammation
      1 hjärnhinneinflammationer
      1 hjärnhinnevätskan
     20 hjärnhinnorna
     14 hjärninfarkt
      1 hjärninfektion
     26 hjärninflammation
      1 hjärninflammationen
      1 hjärnkirurgi
      1 hjärnkomponenter
      1 hjärnlob
      1 hjärnmalaria
      1 hjärnmaterial
      2 hjärnmetastaser
      1 hjärnnhinnorna
      3 hjärnödem
      2 hjärnområden
      1 hjärnoperationer
      7 hjärnor
      1 hjärnparenkym
      1 hjärnparenkymet
      2 hjärnpåverkan
      1 hjärnryggmärgsvätska
      2 hjärnrytmer
      1 hjärnscanning
      1 hjärnscanningsstudier
      2 hjärnsjukdom
      2 hjärnsjukdomar
     17 hjärnskada
      2 hjärnskadade
      3 hjärnskadan
      1 hjärnskaderelaterade
     26 hjärnskador
      1 hjärnskadorna
      1 hjärnskakning
      1 hjärnskakningars
      1 hjärnskanningar
      1 hjärnslag
      2 hjärnstam
     21 hjärnstammen
      1 hjärnstammens
      1 hjärnstamsdöd
      1 hjärnstimulering
      3 hjärnstruktur
      1 hjärnstrukturen
      1 hjärnstrukturer
      2 hjärnstrukturerna
      4 hjärnsubstans
      2 hjärnsubstansen
      1 hjärntillväxten
      1 hjärntrötthet
      1 hjärntrust
     10 hjärntumör
     25 hjärntumörer
      2 hjärntumörerna
      1 hjärntumörfall
      1 hjärntumörföreningen
      1 hjärntumörspatienter
      1 hjärntumörutveckling
      2 hjärntvätt
      1 hjärntvätta
      3 hjärnvågor
      1 hjärnvågsmönster
      1 hjärnvågsstatus
      1 hjärnvattusot
      6 hjärnvävnad
      9 hjärnvävnaden
      1 hjärnventrikeln
     29 hjärt
     32 hjärta
      1 hjärtåkommor
      1 hjärtalungor
      2 hjärtan
      2 hjärtarytmi
      3 hjärtarytmier
      1 hjärtastma
    176 hjärtat
     84 hjärtats
      1 hjärtatsmuskelceller
      1 hjärtattack
      2 hjärtattacker
      1 hjärtaxelns
      1 hjärtbasen
      5 hjärtbesvär
      1 hjärtboken
      3 hjärtcancer
      1 hjärtcellen
      1 hjärtceller
      1 hjärtekrossarfeber
     10 hjärtfel
      1 hjärtflimmer
      1 hjärtformade
      1 hjärtförmak
      9 hjärtfrekvens
      5 hjärtfrekvensen
      1 hjärtfunktionen
      1 hjärthalva
     47 hjärtinfarkt
      2 hjärtinfarkten
      2 hjärtinsufficiens
      1 hjärtkammare
      2 hjärtkärlbiverkningar
      2 hjärtkärlhälsa
      3 hjärtkärlsjukdom
      8 hjärtkärlsjukdomar
      2 hjärtkärlsystemet
      1 hjärtkateter
      1 hjärtkirurgi
      5 hjärtklaffar
      4 hjärtklaffarna
      1 hjärtklaffarnas
      1 hjärtklaffel
      1 hjärtklaffs
      1 hjärtklaffsdegeneration
      1 hjärtklaffsinfektioner
     11 hjärtklappning
      1 hjärtklappningattacker
      1 hjärtklappningsattacker
      1 hjärtklappningsobehag
      1 hjärtkompressioner
      1 hjärtkontrollen
      1 hjärtkranskärlens
      1 hjärtlevande
      3 hjärtljud
      1 hjärtljuden
      1 hjärtlungfonden
      2 hjärtlungmaskin
      4 hjärtlungmaskinen
      1 hjärtlungmaskinens
      1 hjärtlungmaskiner
      1 hjärtlungoperation
      5 hjärtlungräddning
      1 hjärt�lungtransplantation
      1 hjärtmärkningen
      1 hjärtmärkta
      2 hjärtmedicin
      2 hjärtmediciner
      4 hjärtminutvolym
      2 hjärtmissbildningar
      2 hjärtmuskel
      3 hjärtmuskelceller
      2 hjärtmuskelcellerna
      3 hjärtmuskelinflammation
     11 hjärtmuskeln
      1 hjärtmuskelns
      1 hjärtmuskelskada
      1 hjärtmuskelväggen
      1 hjärtmuskler
      2 hjärtmuskulatur
      4 hjärtmuskulaturen
      1 hjärtmuskulaturens
      1 hjärtoperationer
      6 hjärtproblem
      1 hjärtrelaterade
      1 hjärtrubbningar
      4 hjärtrum
      1 hjärtrummen
      1 hjärtrummens
      1 hjärtrusning
      6 hjärtrytm
      2 hjärtrytmen
      1 hjärtrytmrubbning
      3 hjärtrytmrubbningar
      1 hjärtrytmsrubbningar
      2 hjärtsäck
      8 hjärtsäcken
      1 hjärtsäckens
      3 hjärtsäcksinflammation
      1 hjärtsarkom
      1 hjärtsjuka
     12 hjärtsjukdom
     15 hjärtsjukdomar
      1 hjärtsjuke
      1 hjärtskador
      1 hjärtskärande
      9 hjärtslag
      1 hjärtslagen
      1 hjärtslagens
      1 hjärtslagsfrekvens
      1 hjärtslagsfrekvensen
      1 hjärtsonografi
      1 hjärtspecialist
      1 hjärtspecifika
      2 hjärtspetsen
      1 hjärtstatusen
     15 hjärtstillestånd
      1 hjärtstilleståndet
     11 hjärtstopp
      1 hjärtstoppsregistret
     49 hjärtsvikt
      4 hjärtsvikten
      1 hjärtsviktssymptom
      1 hjärtt
      1 hjärttamponad
      5 hjärttransplantation
      1 hjärttumören
      5 hjärttumörer
      1 hjärttumörerna
      2 hjärtväggen
      1 hjärtverksamheten
      1 hjärtverksamhetpuls
      4 hjässa
      3 hjässan
      1 hjertén
      1 hjo
      1 hjord
      1 hjordar
      1 hjorden
      3 hjort
      2 hjortar
      3 hjortdjur
      1 hjortfluga
      1 hjorthornssalt
      1 hjortmärket
      5 hjul
      1 hjulbent
      1 hjulbenta
      6 hjulbenthet
      1 hjulbentheten
      1 hjuldjur
      1 hjulen
      1 hjulet
      1 hkupa
      1 hl
      7 hla
      3 hlaantigen
      1 hlaantigenerna
      1 hladqballelen
      2 hlagen
      1 hlagener
      1 hlagenerna
      1 hlakomplex
      1 hlamolekyl
      1 hlasystemet
      2 hlatest
      6 hlr
      1 hlrrådets
      1 h�lsa
      1 h�morrhoida
      6 hmta
     18 hn
      1 hncn
      1 hno
      2 hnutbrottet
      9 ho
      1 hö
      2 hobby
      1 hobbyändamål
      1 hobbyskyttar
      1 hobbyverksamhet
      2 hobson
      1 hochcoch
      1 [hocho]ch
      1 hocn
      3 hodgkins
      1 hoechst
      1 hofbarnmorskan
      1 hoffberg
      2 hoffer
      2 hoffman
      1 hoffmann
      7 hofmann
      1 hofmanns
      3 höft
      1 höftbenskammen
      1 höftbrott
      5 höften
      2 höftens
      8 höfter
      3 höfterna
      1 höftkammarna
      1 höftledsbyte
      1 höftledsdysplasi
      1 höftmåttet
      1 höftnära
      1 höftprotesoperationer
      1 höftstusskvoten
    355 hög
    196 höga
      1 högaktiv
      2 höganrikat
      1 högättade
      1 högbelastad
      1 högbelastade
      1 högbladen
      1 högdifferentierade
      2 högdos
      1 högdosbehandling
      1 högdosstrålning
      1 högdragenhet
      1 högeffektslaser
     75 höger
      1 högerförmaksförstoring
      2 högerhänta
      1 högerhjärtat
      1 högerkammaren
      1 högerregeln
      1 högersidiga
      3 högersidigt
      3 högertrafikomläggningen
      1 högertrafikversionen
      1 högexplosiva
      1 högfiberkost
      1 högfluortandkräm
      5 högfrekvent
      2 högfrekventa
      5 högfungerande
      2 högg
      1 högglans
      1 höggradiga
      4 höggradigt
      1 höghastighetsborr
      1 höghastighetsborren
      1 höghöjdsbestigningar
      1 höghöjdseffekter
      1 höghöjdslungödem
      1 höghöjdsmedicin
      1 höghöjdsobservatorier
      1 höghöjdsödem
      1 höghöjdssjukdom
      1 höghöjdsträning
      5 höginkomstländer
      1 högintelligenta
      1 högkaloriföda
      1 högkonjunktur
      1 högkostnadsskydd
      2 högkvalitativa
      2 högkvarter
      1 högländerna
      1 höglandet
      1 högläsningen
      1 högläsningsproblem
      1 högljudd
      2 högljutt
      2 högmolekylära
      3 högpresterande
      1 högprioriterade
     34 högra
    265 högre
      1 högrest
      1 högrisk
      1 högriskbeteende
      1 högriskbeteenden
      1 högriskgrupp
      1 högriskgruppen
      3 högriskgrupper
      1 högrisklaboratorium
      1 högrisktyper
      8 högskola
      6 högskolan
      1 högskolebehörighet
      1 högskoleexamen
      1 högskoleförordningen
      1 högskolemässighet
      8 högskolepoäng
      1 högskoleprovet
      4 högskolereformen
      1 högskolestudier
      1 högskoleutbildad
      7 högskoleutbildning
      1 högskoleutbildningar
      1 högskoleutbildningarna
      6 högskoleverket
      1 högskoleverketoch
      3 högskoleverkets
      8 högskolor
      1 högskolorna
      1 högsmittsam
      1 högsommaren
      2 högspänning
      1 högspänningen
      1 högspänningsfält
      2 högspecialiserad
     36 högst
     42 högsta
      1 högstadieskola
      1 högstadiet
      1 högstående
    130 högt
      2 högtalare
      1 högthöga
      1 högtidsuniform
      1 högtrycksmodifikationer
      1 högtrycksstvätt
      1 högupplösande
      1 högvärdigt
      1 högvarv
      1 högväxt
      1 högvuxna
      1 hohenheim
      1 höije
      1 höj
     18 höja
      1 höjas
     39 höjd
      6 höjda
      4 höjden
     13 höjder
      1 höjdes
      1 höjdläget
      3 höjdled
      1 höjdpunkt
     17 höjdsjuka
      1 höjdsjukesymtom
      1 höjdskillnader
      1 höjdssjuka
      9 höjer
      4 höjning
      1 höjningen
     11 höjs
      3 höjt
      1 höjts
      1 holarctica
      1 holbrooki
      1 holdingbolag
      1 holgers
      1 holism
      1 holismen
      3 holistisk
      3 holistiska
      1 holistiskt
      1 höljande
      1 höljd
      4 hölje
      1 höljeförsett
      1 höljeprotein
      2 höljet
      1 höljt
     11 höll
      7 holland
      1 holländare
      1 holländarna
      3 holländska
      1 holländskt
      1 hollerküchle
      1 hollerschöberl
      9 hölls
      1 hollywoods
      1 hollywoodskådespelare
      3 holm
      1 holmes
      1 holmgren
      2 holmiensis
      1 holochlorus
      1 holografiskt
      1 holotyp
      2 hölsterblad
      1 hölsterbladet
      2 homa
      1 homaopatisk
      1 home
      1 homeland
      5 homeopat
      1 homeopaten
      5 homeopater
      1 homeopaterna
      1 homeopathic
      1 homeopathy
     29 homeopati
      1 homeopatiförespråkare
      2 homeopatika
      1 homeopatiker
     17 homeopatin
      3 homeopatins
      4 homeopatisk
     25 homeopatiska
      5 homeopatiskt
      1 homeopatmedel
      1 homeopraktiker
      1 homeos
      7 homeostas
      1 homeostasen
      1 homeostatisk
      1 homeostatiskt
      2 homeros
      1 hominider
      3 hominis
      4 homo
      1 homocysteinemi
      2 homoeopathic
      1 homoeroticism
      1 homofon
      1 homofoner
      1 homogen
      1 homogena
      1 homogeniserad
      1 homolog
      1 homonet
      1 homonym
      1 homosexualitet
      1 homosexuell
     16 homosexuella
      1 homotoxicosis
      1 homotoxikologi
      1 homotoxikos
      3 homozygot
      1 homozygota
      1 homunculi
    141 hon
      6 hona
      1 höna
     26 honan
      5 honans
      4 honblommor
      1 honblommorna
      1 honblommornas
      2 hondjur
      1 honeymoon
      1 hong
      1 hongamofyten
      2 hongkong
      2 hongkonginfluensan
      3 honhan
      1 honkotten
      1 honkottenbäret
      2 honlig
      3 honliga
      1 honmasken
     33 honom
      2 honomhenne
     31 honor
      2 honorganet
     13 honorna
      2 honornas
      1 honplantan
      2 höns
      2 hönsabane
      2 hönsägg
      1 hönsfåglar
      1 hönsfjädrar
      1 honsporangiets
      8 honung
      1 honungs
      1 honungspung
      2 honungsskivling
      5 honungsskivlingar
      3 honungsskivlingarna
      5 honungsskivlingen
      4 honungsskivlingens
      1 honungsskivlingsarten
      1 honvaraner
      1 höök
      1 hookeri
      2 hoorn
      1 hoover
      1 hopade
      1 hopböjd
      1 hopdragningar
      1 hopen
      2 hopfogad
      2 hopkins
      1 hopklämning
     13 hopp
      5 hoppa
      2 hoppades
      1 hoppande
      3 hoppar
      3 hoppas
      1 hoppat
      2 hoppfullhet
      1 hoppingivande
      2 hoppkräftan
      5 hoppkräftor
      2 hoppkräftorna
      2 hopplösa
      5 hopplöshet
      1 hopplöst
      1 hoppträning
      1 hopsnurrade
      1 hoptrasslad
      1 hoptryckt
      1 hopvikt
     26 hor
    130 hör
      2 hora
     25 höra
      6 hörande
      7 hörapparat
      2 hörapparaten
      1 hörapparatenhörsnäcka
      4 hörapparater
      1 hörapparaterna
      5 höras
      2 hörbara
      1 hörbarhet
      1 hörbarhetsområde
      1 hörcentral
     10 hörde
      1 hordein
      1 hordeiner
      1 hörhjälpmedel
      1 horisontala
      1 horisontalis
      1 horisontalstammen
      9 horisontell
      5 horisontella
      8 horisontellt
      2 horisonten
      2 horizon
      1 horkarl
      1 hörlur
      2 hörlurar
      1 hormesis
     87 hormon
      1 hormonaktivitet
      2 hormonaktiviteten
      2 hormonbalansen
      1 hormonbaserade
      9 hormonbehandling
      2 hormonbehandlingar
      1 hormonblockerande
      1 hormoncykel
      1 hormone
     10 hormonell
     17 hormonella
      3 hormonellt
    124 hormoner
     45 hormonerna
      3 hormonernas
      1 hormoners
     46 hormonet
      1 hormonfluktuationer
      3 hormonförändringar
      1 hormonfrisättande
      1 hormongrupper
      1 hormonhalten
      1 hormonhalter
      1 hormoniellt
      1 hormoninsöndring
      1 hormoninsöndringen
      1 hormoninverkan
      1 hormonkoncentrationer
      1 hormonkörtel
      5 hormonkörtlar
      1 hormonkörtlarna
      1 hormonläkemedel
      1 hormonlika
      2 hormonliknande
      1 hormonmängden
      1 hormonmodulerare
      1 hormonnedbrytningsprodukt
      1 hormonnivå
      6 hormonnivåer
      8 hormonnivåerna
      3 hormonnivån
      1 hormonöverkänslighet
      1 hormonplåster
      1 hormonpreparat
      6 hormonproducerande
      3 hormonproduktion
      5 hormonproduktionen
      1 hormonprofil
      1 hormonprover
      1 hormonresponselement
      6 hormonrubbningar
      2 hormonspiral
      1 hormonspiraler
      2 hormonstörande
      1 hormonstörning
      1 hormonstörningar
      2 hormonsvängningar
      2 hormonsystem
      1 hormontabletter
      2 hormonvärden
      1 hormoslyr
      7 horn
      4 hörn
      1 hornblände
      2 horne
      1 hörnen
      2 horners
      3 hornet
      2 hörnet
      1 hornets
      1 hornhinna
     10 hornhinnan
      1 hornhinnans
      2 hornhinnor
      1 hornlager
      1 hornlagret
      1 hornråg
      1 hörntänderna
      3 horridum
      2 hörs
      1 hörsammar
      3 horsbrott
      3 horsbrottet
      1 horsehoof
     28 hörsel
      2 hörselbenen
      1 hörselbortfall
      1 hörselcentrum
      1 hörselförändringen
      1 hörselförlust
      2 hörselgångarna
      3 hörselgången
      4 hörselhallucination
      1 hörselhallucinationen
     11 hörselhallucinationer
      3 hörselhallucinationerna
      1 hörselkliniken
      1 hörselläkare
      9 hörseln
     22 hörselnedsättning
      3 hörselnedsättningar
      3 hörselnedsättningen
      1 hörselnedsättninghörselskador
      1 hörselnerv
      5 hörselnerven
      1 hörselnerverna
      1 hörselnervsinflammation
      1 hörselns
      1 hörselrest
      1 hörselrester
      1 hörselsinne
      5 hörselskada
      6 hörselskadade
      1 hörselskadadedöva
      1 hörselskadades
      2 hörselskador
      1 hörselskydd
      1 hörselskyddhörselproppar
      1 hörselslingateleslinga
      1 hörselsnäcka
      7 hörselsnäckan
      1 hörselsystem
      1 hörseltekniska
      3 hörseltest
      3 hörselundersökningar
      1 hörselupplevelsen
      1 hörselvården
      1 hörselvårdsutredningen
      1 hörslang
      1 hörsneloka
      3 hört
      1 hörtelefon
      2 hörtröskel
      2 hörtröskeln
      1 hörupplevelse
      1 hörupplevelserna
   1742 hos
      1 hosack
      1 hosmän
      4 hösnuva
      1 hösnuvesymtom
      1 hospisvård
     12 hospital
      3 höst
     69 hosta
      2 höstadonis
      7 hostan
      6 hostar
      4 hostas
      1 hostat
      3 hostattackerna
      1 höstblåsor
      2 hostdämpande
     27 hösten
      1 höstenvintern
      1 hosthäva
      5 hostmedicin
      1 hostmedicinen
      2 hostmediciner
      1 hostning
      2 hostningar
      1 hostningen
      1 hostreflexen
      1 hostretande
      1 höstsås
      1 höstterminen
     45 hot
      3 hota
     10 hotad
      3 hotade
      2 hotande
      4 hotar
      4 hotas
      1 hotat
      1 hotel
      1 hotell
      1 hotellbranschen
      1 hoten
      3 hotet
      1 hotfull
      8 hotfulla
      1 houghton
      1 hounsfield
      1 hour
      6 house
      1 houses
      1 houston
      1 houyhnhnm
      2 hov
      1 hovbarnmorskan
      1 hovdjur
      1 hovdjuren
      1 hovgräs
      1 hovrätt
      1 hovtångliknande
      3 howard
      1 hoxd
      1 hoysala
      6 hp
      3 hpaaxeln
      1 hpaaxelns
      1 hparametrar
      1 h�pital
      1 h�pnos
      1 h�pochóndrios
      2 hppd
     12 hpv
      1 hpvviruset
      2 h�r
      1 hre
      1 hreceptorblockerare
      1 hridaya
      2 hrt
      2 hrv
      1 hsan
      1 hsiung
      3 hsl
      4 hso
      3 hsp
      1 hsv
      2 hta
      1 h�tel
      1 htlvi
      2 htlviii
      3 htt
      1 httpdrgabormatecom
      1 httpenwikipediaorgwikianthrax
      1 httpflickansaarabloggse
      1 httpreliefwebintdisasterepslv
      1 httpsratseyrkenperfusionist
      1 httpswwwfacebookcomgroups
      1 httpswwwhavochvattensehavfiskefritidfritidsbatarrenbatbottenhtml
      1 httpswwwncbinlmnihgovpmcarticlespmcncbisevere
      1 httpswwwyoutubecomchannelucfxrjlxtzqodkjiyawvideos
      1 httpwwwaftonbladetsekropphalsaarticleabserviceprint
      1 httpwwwakademiskasesvverksamheterneurokirurgi
      1 httpwwwastmaoallergiforbundetse
      1 httpwwwcholangiocarcinomaorg
      1 httpwwwdnsenyhetersvarareattfaljusterapi
      1 httpwwwdukoralse
      1 httpwwwdyslexiorg
      1 httpwwwfdbnu
      1 httpwwwhealthcommunitiescomurologiskaakutfallpriapismshtml
      1 httpwwwkarolinskaseverksamheternasklinikerenheterneurokirurgiskakliniken
      1 httpwwwkarolinskaseverksamheternasklinikerenheterneurokirurgiskaklinikenforskninginomneurokirurgi
      1 httpwwwkarolinskaseverksamheternasklinikerenheterneurokirurgiskaklinikenfunktionellneurokirurgi
      1 httpwwwlakartidningenseenginephparticleid
      1 httpwwwlakartidningensefunctionsoldarticleviewaspxarticleid
      1 httpwwwlioseomlandstingetverksamhetersinnescentrumneurokirurgiskaklinikenilinkoping
      1 httpwwwmedluseklinvetlundneurokirurgi
      4 httpwwwncbinlmnihgovpubmed
      1 httpwwwncbinlmnihgovpubmedncbi
      1 httpwwwncbinlmnihgovpubmedncbihigh
      1 httpwwwneuropharmumuseominstitutionenenheterklinneurovet
      1 httpwwwneurouuseresearchneurosurgerylanguageid
      1 httpwwwnewsmedicalnethealthsymptomsofcyanosisswedishaspx
      1 httpwwwrcorg
      1 httpwwwsahlgrenskasesvsuvardhygien
      1 httpwwwsciencedirectcomsciencearticlepiisscience
      1 httpwwwslusesvomslufristaendesidoraktuelltallanyheternyametoderfordiagnosavvingelsjukahoskatt
      1 httpwwwsmittskyddsinstitutetsesjukdomarmjaltbrand
      1 httpwwwsocialstyrelsenseovanligadiagnoserklippeltrenaunayssyndrom
      1 httpwwwsvenskaktsnatverketse
      1 httpwwwsvtsenyhetervetenskapjaktenpasmittansursprung
      1 httpwwwtandlakartidningensemediapdf
      1 httpwwwtopfholocaustde
      1 httpwwwvardguidensesjukdomarochradomradensjukdomarochbesvarmjaltbrand
      1 httpwwwwebfinansercomnyheterid
      1 httpwwwwhointwerwerenindexhtml
      1 hu
      1 hua
      1 hubel
    108 hud
      2 hudabscesser
      1 hudåkomma
      1 hudåkommor
      1 hudallergitester
      1 hudar
      1 hudavfall
      1 hudavlagringar
      3 hudbakterier
      2 hudbarriären
      1 hudbesvär
      2 hudbiopsi
      1 hudbitar
      1 hudbitarna
      1 hudblödningar
     18 hudcancer
      1 hudcancerpatienten
      2 hudceller
      2 huddesinfektion
      4 huddinge
    306 huden
     20 hudens
      1 hudepitel
      2 hudfärg
      1 hudfärgad
      1 hudfärgade
      2 hudfärgat
      1 hudfläcken
      1 hudflagor
      1 hudflik
      1 hudflikar
      1 hudförändring
      6 hudförändringar
      2 hudförtunning
      1 hudgenomblödningen
      1 hudimplantat
      1 hudinfektion
     11 hudinfektioner
      3 hudinflammation
      2 hudinflammationer
      2 hudirritation
      1 hudkänseln
      1 hudkänslighet
      1 hudklinik
      1 hudkliniker
      5 hudkontakt
      1 hudkörtel
      5 hudkräm
      1 hudkrämen
      6 hudkrämer
      3 hudlager
      2 hudlagren
      5 hudlagret
      1 hudläkare
      1 hudlesion
      1 hudlesioner
      2 hudlotion
      1 hudmothudkontakt
      1 hudoch
      1 hudödem
      2 hudområde
      3 hudområden
      1 hudområdet
      1 hudömsning
      1 hudpartier
      1 hudporfyrierna
      2 hudprover
      1 hudpsoriasis
      1 hudreaktion
      1 hudreaktioner
      1 hudrispa
      3 hudrodnad
      1 hudrodnaden
      1 hudrodnader
      4 hudsår
      4 hudsjukdom
      7 hudsjukdomar
      2 hudsjukdomen
      1 hudskada
      3 hudskador
      1 hudskick
      1 hudson
      1 hudspecialist
      1 hudsträng
      1 hudsträngen
      1 hudsvamp
      1 hudsvampinfektion
      1 hudsvullnaderna
      1 hudsymptomen
      4 hudsymtom
      1 hudtemperatur
      1 hudtest
      1 hudtester
      2 hudtonen
      1 hudtransplantion
      1 hudtuberkulos
      1 hudtumör
     12 hudutslag
      1 hudvalk
      1 hudvalkar
      1 hudvård
      2 hudvårdsprodukter
      1 hudvävnad
      6 hudytan
      2 huehuetenango
      1 hufvudena
      1 hugg
      3 hugga
      1 hugger
      1 huggkänslor
      2 huggorm
      2 huggormar
      1 huggormen
      1 huggsår
      1 huggtand
      4 huggtänder
      1 huggtänderna
      2 hughes
      1 hughlings
      1 hugo
      1 huitlacoche
      1 hukande
      2 hullingar
      1 hullingförsedd
      1 humalog
     13 human
     10 humana
      3 humanbiologi
      1 humanceller
      1 humanfall
      1 humanfallen
      1 humanfysiologin
      1 humani
      2 humaniora
      1 humanist
      2 humanistisk
      7 humanistiska
      1 humanitära
      1 humankapital
      1 humanmedicin
      1 humanmedicinen
      1 humanpatogen
      1 humanpatogena
      1 humans
     17 humant
      1 humbled
      1 humboldt
      1 humen
      1 humerus
      1 humilis
      1 humira
      1 humla
      1 humle
      1 humlor
      2 humor
      5 humör
      2 humoral
      3 humorala
      4 humoralpatologi
      5 humoralpatologin
      1 humoralpatologiska
      4 humöret
      1 humoristiska
      1 humoristiskt
      1 humörstörningar
      1 humörsvängingarsvårighet
     12 humörsvängningar
      1 humphrey
      4 humphry
      1 humrar
     34 hund
     61 hundar
      5 hundarna
      2 hundbett
      1 hunddagis
     31 hunden
      4 hundens
      1 hundetjenster
      1 hundförsäkringen
      2 hundhybrid
      1 hundliv
      1 hundloka
     27 hundra
      1 hundraårskriget
      2 hundrade
      1 hundraprocentig
      2 hundraser
      1 hundrastgårdar
      2 hundratal
      1 hundratalas
     11 hundratals
      1 hundratusen
      4 hundratusentals
      1 hundred
      6 hundrova
      1 hundrovesläktet
      1 hundrovor
      1 hundsjukdomar
      1 hundteamet
      1 hundtjänst
      1 hundvalpar
     14 hunger
      2 hungerdämpande
      2 hungerkänslor
      2 hungerkänslorna
      3 hungern
      1 hungerscentrum
      5 hungersnöd
      1 hungersnöden
      5 hungrig
      5 hungriga
      1 hunnen
     11 hunnit
      1 hunt
      1 hunter
      5 huntingtin
      5 huntingtons
      1 hunza
      1 huor
    569 hur
      1 hurme
      1 hurudana
     71 huruvida
     15 hus
      1 husägare
      1 husandar
      1 husarbete
      1 husbränder
      1 husdamm
      2 husdammskvalster
     14 husdjur
      1 husdjurs
      1 husdjursavel
      4 huset
      1 husets
      1 husförhörslängd
      1 husförhörslängden
      3 husgeråd
      2 husgolv
      4 hushåll
      2 hushållen
      2 hushållet
      1 hushållets
      1 hushållning
      1 hushålls
      1 hushållsarbete
      1 hushållsarbetet
      3 hushållsbruk
      1 hushållsdammsugare
      1 hushållshandskar
      1 hushållsmiljö
      2 hushållsnära
      9 hushållspapper
      1 hushållspapperet
      1 hushållssopornabrännbart
      1 hushållssvamp
      1 hushållssysslorna
      1 hushållstrupper
      1 hushållstvål
      1 hushållstvätten
      2 huskur
      2 huskurer
      1 huskvarna
      1 husläkar
      1 husläkare
      1 husläkarmottagning
      1 husmanskost
      1 husmusens
      1 husockupation
      2 husrannsakan
      1 husrannsakningsorder
      1 huss
      1 husse
      1 husserl
      9 hustru
      3 hustrun
      1 hustrur
      1 hustrurs
      1 husvagnsekipage
      2 hutchinson
      6 hutchinsongilfords
      1 huvdkontor
     43 huvud
      1 huvudakligen
      3 huvudämne
      1 huvudänden
      1 huvudansvaret
      1 huvudargumentet
      2 huvudartikel
      1 huvudbeståndsdelen
      1 huvudbonad
      1 huvudbonader
      1 huvudbry
      1 huvudceller
      1 huvudcenter
      1 huvuddel
      3 huvuddelar
      1 huvuddelarna
     11 huvuddelen
      2 huvuddrog
      1 huvuddrogen
      3 huvuden
     69 huvudet
      5 huvudets
      1 huvudfaktor
      1 huvudfårans
      1 huvudförfattaren
      2 huvudfunktionen
      1 huvudgrenar
      5 huvudgrupper
      3 huvudgrupperna
      1 huvudhår
      1 huvudhöjd
      1 huvudingrediens
      1 huvudinriktning
      1 huvudkanal
      1 huvudkaraktären
      1 huvudkategori
      1 huvudkategorier
      1 huvudkedjan
      3 huvudklasser
      1 huvudklassificeringar
      1 huvudkomponenter
      1 huvudkomponenterna
      8 huvudkontor
      2 huvudkontoret
      1 huvudkriterier
      1 huvudkriterierna
      1 huvudkrona
      1 huvudled
      3 huvudleden
      1 huvudlinjer
      2 huvudlöss
      1 huvudlusen
      2 huvudlusens
      2 huvudman
      1 huvudmannaskap
      1 huvudmannaskapet
      3 huvudmannen
      1 huvudmetaboliten
      1 huvudmissbruket
      1 huvudnamnet
      1 huvudnyckel
      1 huvudomfång
      1 huvudområden
      1 huvudorsak
      5 huvudorsaken
      1 huvudort
      1 huvudorten
      1 huvudperson
      7 huvudpersonen
      3 huvudpersoner
      1 huvudposition
      1 huvudprincip
      1 huvudprincipen
      1 huvudprinciper
      1 huvudpulsådern
      1 huvudregionen
      2 huvudriktningar
      1 huvudrollerna
      1 huvudrollsinnehavarens
      1 huvudrörelse
      2 huvudrörelser
      1 huvudrot
     32 huvudsak
      3 huvudsaklig
     64 huvudsakliga
      1 huvudsaklige
    100 huvudsakligen
      1 huvudsaksigen
      1 huvudsatser
      1 huvudsjukdomen
      2 huvudskada
      1 huvudskål
      1 huvudskålens
      1 huvudskälet
      1 huvudspänningen
      1 huvudstäder
      1 huvudställningar
      1 huvudställningskomfort
      2 huvudstammen
      1 huvudstammens
      2 huvudsyfte
      1 huvudsymptom
      3 huvudsymtom
      1 huvudtecken
      1 huvudtema
      1 huvudteorier
      1 huvudtillverkaren
      7 huvudtyper
      1 huvudtyperna
      2 huvuduppgift
      1 huvudvägen
      1 huvudvärden
    106 huvudvärk
      5 huvudvärken
      3 huvudvärksdiagnos
      2 huvudvärksformer
      1 huvudvärksformerna
      1 huvudvärkssjukdomar
      1 huvudvärkssjukdomarna
      1 huvudvärksspecialister
      1 huvudväxel
      1 huvudverktygen
      1 huxley
      1 huxtable
      1 hvor
      1 hwad
      1 hwarang
      1 hwarest
     10 hy
      1 hyacintväxter
      1 hyalint
      1 hyalinum
      1 hyaloidea
      1 hyaluronidas
      4 hyaluronsyra
      4 hybrid
      1 hybrida
      1 hybridcellen
      1 hybriden
      5 hybrider
      1 hybridgullregn
      1 hybridisera
      2 hybridom
      1 hybridomceller
      1 hybridomer
      2 hybridomteknologi
      1 hybridomteknologin
      1 hybridteknik
      1 hydatidos
      1 hydatitosa
      1 hyde
      1 hydōr
      1 hydrargentum
      1 hydrargyros
      1 hydrater
      1 hydration
      5 hydratisering
      1 hydraulvätska
      1 hydrering
      1 hydrid
      1 hydroargentum
      1 hydrocarbon
      7 hydrocefalus
      5 hydrocephalus
      3 hydrofil
      4 hydrofila
      2 hydrofilt
      2 hydrofob
      6 hydrofoba
      2 hydrofobi
      2 hydrofobt
      1 hydrofon
      1 hydrogeneras
      1 hydrokephalos
      6 hydrokinon
      1 hydrokloridformen
      2 hydrokortison
      5 hydrolys
      2 hydrolysen
      1 hydrolysera
      2 hydrolyserar
      1 hydrolyseras
      1 hydromorfon
      5 hydronefros
      1 hydronium
      1 hydroöstron
      1 hydrophids
      3 hydror
      5 hydrostatiska
      1 hydrostatiskt
      1 hydroterapi
      1 hydroxi
      1 hydroxiandrostenon
      3 hydroxiantracen
      1 hydroxiantracenderivat
      1 hydroxiapatit
      1 hydroxibensoesyra
      1 hydroxicyklohexadienon
      1 hydroxid
      1 hydroxiderivatet
      1 hydroxidjoner
      1 hydroxietylstärkelse
      1 hydroxifenol
      3 hydroxigrupp
      2 hydroxigruppen
      2 hydroxigrupper
      1 hydroxiketoner
      2 hydroxiprogesteron
      1 �hydroxiprogesteron
      1 hydroxipropansyra
      1 hydroxisyror
      1 hydroxyecdysteron
      1 hydroxyindolacetat
      3 hydroxylapatit
      3 hydroxylation
      1 hydroxylera
      1 hydroxyleras
      1 hydroxylering
      1 hydroxylerna
      4 hydroxylgrupp
      4 hydroxylgruppen
      4 hydroxylgrupper
      1 hydroxyljoner
      1 hydroxylradikaler
      1 hydrozoer
      2 hyemalis
      1 hyena
      3 hyfer
      3 hyferna
      1 hyfgrenar
      1 hyfsat
      1 hyggen
      3 hygieia
     39 hygien
      1 hygienartikel
      1 hygienartikels
      5 hygienartiklar
      1 hygiene
      3 hygienen
      2 hygienens
      1 hygienföreskrifterna
      2 hygienisk
     11 hygieniska
      1 hygieniskdietetiska
      1 hygieniskdietisk
      3 hygieniskt
      1 hygiennivån
      1 hygienområdet
      1 hygienpraxis
      1 hygienproblem
      1 hygienprodukt
      7 hygienprodukter
      1 hygienregler
      1 hygienrutiner
      1 hygientekniker
      1 hygienvanan
      1 hygrophilus
      1 hygroskopisk
      1 hygroskopiskt
      1 hylander
      1 hylden
      1 hyll
      1 hylla
      1 hyllade
      1 hyllades
      2 hyllar
      2 hylle
      4 hylleblad
      2 hyllebladen
      1 hyllebuske
      1 hyllerester
      1 hyllesaft
      1 hyllningar
      1 hyllningsgala
      1 hyllor
      1 hylsan
      1 hylsor
      1 hymenium
      1 hymenochaetaceae
      1 hymenoptera
      1 hyn
      1 hyoglossus
      1 hyoidbenet
      5 hyoscyamin
      1 hyoscyamus
      2 hyper
      1 hyperactiveimpulsive
      1 hyperactivity
     15 hyperacusis
      1 hyperacusisljudöverkänslighet
      1 hyperaktiv
      2 hyperaktiva
     14 hyperaktivitet
      2 hyperaktivitetimpulsivitet
      1 hyperaktivitetsstörningar
      1 hyperaktivt
     15 hyperakusi
     11 hyperalgesi
      3 hyperammonemi
     13 hyperandrogenism
      1 hyperandrogenismen
      1 hyperandronenism
      1 hyperbar
      1 hyperbarmedicin
      3 hyperbilirubinemi
      1 hypercapnia
      2 hyperemotionella
      1 hyperestesi
      1 hyperexhalterad
      1 hyperfagi
      1 hyperfiltrerar
      4 hyperfunktion
      2 hyperglykemi
      2 hyperglykemiskt
      1 hypergonadism
      2 hypergonadotropism
      4 hypergrafi
     11 hyperhidros
      1 hyperhidrosis
      1 hyperhörsel
      1 hyperinflation
      1 hyperinsulinemi
      1 hyperinsulinism
      6 hyperkalcemi
      4 hyperkalemi
      1 hyperkalemin
      2 hyperkapni
      9 hyperkeratos
      1 hyperkeratosen
      1 hyperkeratotiskt
      1 hyperkinesi
      1 hyperkinetic
      1 hyperkinetisk
      7 hyperkolesterolemi
      4 hyperkortisolism
      1 hyperlexi
      1 hypermenorré
      1 hypermobil
      2 hypermobilitet
      1 hyperosmolärt
      3 hyperöstrogenism
      1 hyperparatyreos
      1 hyperpigmenterad
      1 hyperpigmenterat
      3 hyperpigmentering
      5 hyperplasi
      1 hyperplasier
      2 hyperplastisk
      1 hyperplastiskt
      1 hyperpolariserat
      1 hyperpolariseringen
      1 hyperproduktion
     10 hyperprolaktinemi
      6 hyperreaktivitet
      1 hyperreflexi
      1 hypersekretion
      1 hypersensitiviten
     16 hypersensitivitet
      1 hypersensitivitetsreaktion
     17 hypersomni
      1 hypersomnier
      1 hypersomnin
      1 hyperstimulering
      4 hypertelorism
      1 hypertelorismen
      4 hypertension
      3 hypertermi
      1 hyperthyreos
      2 hyperton
     10 hypertoni
      3 hypertriglyceridemi
     10 hypertrofi
      1 hypertrofiskcellvävnads
      2 hypertymesi
      1 hypertymestisk
      1 hypertymestiskt
      3 hypertyreos
      1 hypertyroidism
      1 hyperuppblåsta
      6 hyperurikemi
     15 hyperventilation
      2 hyperventilationen
      2 hyperventilera
      1 hyperventilerar
      1 hyperventilering
      1 hyperventileringen
      1 hyperviskositet
      1 hyperviskositetssymtom
      4 hypestesi
      1 hypestesin
      1 hypestisti
      1 hyphodontia
      2 hypnagog
      3 hypnagoga
      1 hypnogramdormogram
      2 hypnopomp
      2 hypnopompa
     24 hypnos
      1 hypnosens
      1 hypnotiserad
      3 hypnotiserade
      2 hypnotisk
      9 hypnotiska
      1 hypnotiskt
      4 hypnotisören
      1 hypnotisörens
      1 hypo
      1 hypoaktiv
      1 hypoaktivitet
      1 hypoalbuminemi
      1 hypoallergeniska
      3 hypoandrogenism
      1 hypochlorous
      2 hypoderma
      1 hypoemotionalitet
      1 hypoestrogenism
      1 hypoestrogenismen
      1 hypofarynx
      2 hypofys
      1 hypofysadenom
      3 hypofysär
     57 hypofysen
     14 hypofysens
      1 hypofysfunktion
      1 hypofyshämmande
      1 hypofyshormon
      1 hypofyshormoner
      5 hypofysinsufficiens
      1 hypofysiotropa
      2 hypofysområdet
      1 hypofystumör
      1 hypofystumören
      5 hypofystumörer
      1 hypogeusi
      1 hypoglossus
     13 hypoglykemi
      4 hypoglykemisk
     12 hypogonadism
      1 hypogonadotrop
      4 hypogonadotropism
      4 hypokalcemi
      1 hypokalcemiska
      7 hypokalemi
      1 hypokinesi
      1 hypokinetisk
      2 hypoklorit
      2 hypokloriter
      3 hypokloritsyra
      1 hypoklorsyra
     13 hypokondri
      2 hypokondriker
      2 hypokondrin
      1 hypokondrium
      1 hypokretin
      1 hypokrom
     21 hyponatremi
      5 hypoöstrogenism
      1 hypoparathyreoidism
      1 hypopharynx
      1 hypopigmenterade
      1 hypopigmenterat
      1 hypopituitarism
      1 hypopiuitarism
      1 hypopnéer
      1 hypopolarisering
      1 hypopyon
      7 hyposensibilisering
      4 hyposensitivitet
      5 hypospadi
      1 hyposplenism
     40 hypotalamus
      1 hypotalamushypofyskönskörtelsystemet
     11 hypotermi
     28 hypotes
     15 hypotesen
     12 hypoteser
      1 hypoteserna
      1 hypotesprövning
      1 hypotetisk
      1 hypotetiska
     16 hypothalamus
      1 hypothesis
      1 hypoton
      3 hypotoni
     22 hypotyreos
      1 hypotyroida
      3 hypotyroidism
      1 hypotyroidliknande
      2 hypoventilation
      6 hypovolemi
      1 hypovolemisk
      4 hypoxemi
     17 hypoxi
      1 hypoxin
      1 hypoxisk
      1 hypsignathus
      1 hyra
      1 hyrbröder
      1 hyresgäst
      1 hyresgästen
      1 hyreshus
      2 hyresrätt
      1 hyresrätten
      2 hyresvärden
      1 hyrocefalus
      1 hyrs
      1 hyrsyskon
      1 hyrsystrar
      1 hysa
      5 hyser
      2 hyskor
      1 hystera
      3 hysterektomi
     16 hysteri
      1 hysteria
      1 hysterikor
      2 hysterin
      1 hysteripatienter
      5 hysterisk
      6 hysteriska
      1 hysteroskop
      3 hysteroskopi
      1 hyvac
     23 hz
  18683 i
      1 [i
      1 ia
      1 iaea
      1 iaeas
      4 iaktta
      1 iakttaga
      1 iakttagande
      1 iakttagandet
      1 iakttagbara
      2 iakttagelse
      3 iakttagelser
      4 iakttagits
      2 iakttar
      5 iakttas
      1 iakttog
      2 iakttogs
      1 ian
      1 iands
      1 iarc
      1 iast
      1 iasttransliteration
      1 iatraléiptai
      1 iatrogen
      2 iatrogena
      1 iband
      1 ibererna
      1 iberisk
    572 ibland
      1 iblandade
      1 ibm
      1 iboga
      1 ibogain
      1 ibot
      1 ibotensyra
      2 ibs
      1 ibsa
      1 ibsen
      5 ibuprofen
      3 ica
      1 icamreceptorer
      1 icchp
     90 icd
      2 icdcm
      1 icds
      1 icdse
      1 iceller
      1 icer
      1 ichimura
      1 ickaadministrativt
     57 icke
      2 ickeakuta
      2 ickeallergisk
      1 ickeallvarlig
      2 ickeanimalisk
      1 ickeariskt
      1 ickeatman
      1 ickeavvikare
      1 ickebakteriell
      1 ickebakteriella
      1 ickebestrålade
      1 ickebleknande
      2 ickebrännbar
      1 ickebrustet
      1 ickecellulär
      1 ickedömande
      2 ickeendemiska
      1 ickeenzymatisk
      1 ickeenzymatiska
      1 ickeepileptiker
      2 ickeexisterande
      1 ickeexplosiva
      1 ickefalsifierbar
      4 ickefarmakologisk
      1 ickefientliga
      1 ickeflytande
      1 ickeformell
      1 ickeförvärvsarbetande
      1 ickefotosyntetiserande
      1 ickefruktbärande
      1 ickefysiologisk
      1 ickegiftiga
      2 ickegravida
      1 ickehemolytiska
      1 ickehereditära
      1 ickehumana
      2 ickeimmun
      1 ickeimmuna
      1 ickeimmunförmedlade
      1 ickeimmunologisk
      3 ickeinfektiös
      3 ickeinfektiösa
      1 ickeinsulinkrävande
      6 ickeinvasiv
      2 ickeinvasiva
      1 ickejoniserande
      1 ickekirurgisk
      2 ickekirurgiska
      1 ickekliande
      1 ickekliniska
      1 ickekodande
      1 ickekonstruktiva
      3 ickekriminella
      2 ickekriminellt
      1 ickekroppslig
      1 ickekroppsliga
      1 ickekvantitativa
      1 ickemanifesterad
      2 ickemänniskoapor
      4 ickemedicinska
      2 ickemedicinskbehandling
      1 ickemedicinskt
      1 ickemelankoliska
      1 ickemelanom
      1 ickemetalliskt
      1 ickemilitära
      1 ickemineraliserad
      1 ickemonetär
      2 ickenaturlig
      2 ickeneurogena
      1 ickenormal
      1 ickenormala
      1 ickenukleosid
      1 ickeoperativ
      1 ickeorganisk
      1 ickeortogonala
      1 ickeparasitiska
      1 ickeproteinbundna
      1 ickepsykopatisk
      1 ickeradioaktiv
      1 ickeradioaktiva
      1 ickereaktiva
      2 ickeremsömn
      1 ickeresistent
      1 ickeresistenta
     10 ickerökare
      1 ickerörliga
      1 ickesexuellt
      1 ickesjukdom
      6 ickesmåcelliga
      1 ickespecialiserade
      3 ickespecifik
      2 ickespecifika
      1 ickespråklig
      2 ickespråkliga
      1 ickespridd
      1 ickestandardiserad
      1 ickestatliga
      4 ickesteroida
      1 icketoxiska
      1 icketraumatiska
      2 ickeundvikandeterapi
      1 ickeupplysta
      1 ickevaccinerade
      3 ickevästerländska
      1 ickeverbal
      1 ickeverbala
      1 icnirp
      1 icnirps
      2 icoh
      1 icrp
      4 icsd
      1 icsdkriterierna
      1 id
      4 ida
    308 idag
      1 idarubicin
      5 idé
      8 ideal
      1 ideala
      1 idealiserad
      2 idealiserade
      3 idealisk
      2 idealiska
      3 idealiskt
      1 idealism
      1 idealismen
      1 idealistisk
      1 idealplagg
      4 idealt
      1 idealvikt
      1 ideation
      1 ideatorisk
      1 idédrama
      1 ideell
      3 ideella
      1 ideellt
     17 idéer
      2 idéerna
      1 idéflykt
      1 idégivaren
     17 idegran
      1 idegranars
      1 idegranarten
      9 idegranen
      1 idegranens
      1 idegranplantor
      1 idegransbast
      1 idegransbeståndet
      1 idegransöarna
      1 idegransrunan
      1 idéhistorikern
      1 idéhistoriska
      1 idéhistoriskt
     22 idén
     51 identifiera
      1 identifierad
      8 identifierade
     10 identifierades
      7 identifierar
      9 identifieras
      7 identifierat
      5 identifierats
      8 identifiering
      5 identifikation
      2 identifikationen
      1 identifikatorer
      4 identisk
     10 identiska
      4 identiskt
     12 identitet
      1 identiteten
      1 identitetsskapande
      2 identitetsstörning
      1 identity
      2 ideologi
      3 ideologisk
      2 ideologiska
      2 ideologiskt
      8 ideomotorisk
      1 idiabetes
     10 idiopatisk
      2 idiopatiska
      2 idios
      2 idiosynkrasi
      1 idiosynkrasia
      7 idiot
      2 idiotanstalten
      1 idiotanstalter
      1 idiotbegreppet
      6 idioter
      1 idioterna
      1 idiotes
      6 idioti
      1 idiotundervisning
     12 idisslare
      1 idogt
      1 idol
      1 idoler
      3 idrott
      2 idrottande
      1 idrottandet
      1 idrottar
      3 idrottare
      2 idrottaren
      3 idrotten
      1 idrottens
      2 idrotter
      1 idrottsböcker
      1 idrottsgren
      2 idrottshjärta
      2 idrottskvinnor
      4 idrottsmän
      1 idrottsmassage
      3 idrottsmedicin
      2 idrottsmedicinen
      1 idrottsmekanik
      1 idrottsplatser
      1 idrottspsykologi
      1 idrottsrelaterad
      1 idrottsrelaterade
      2 idrottsskada
      7 idrottsskador
      1 idrottstävlingar
      1 idrottsutövare
      1 idrottsvärlden
      1 idsa
      1 idylliska
      1 ie
      1 iec
      2 ieee
      1 iekg
      1 if
     10 ifall
      1 iförd
      1 ifosfamid
     28 ifråga
     12 ifrågasatt
      1 ifrågasatta
      7 ifrågasätta
      1 ifrågasättande
      1 ifrågasättandet
      5 ifrågasättas
      1 ifrågasätter
      1 ifrågasattes
      6 ifrågasatts
      4 ifrågasätts
     80 ifrån
      1 ifred
      1 ifvitaminbkomplex
      1 ig
      4 iga
      1 iganefrit
     42 igång
      1 igångsatta
      1 igatyp
      7 ige
      2 igeantikroppar
      1 ige�antikroppar
      1 igeantikropparna
      1 igeantikroppsaktivering
      3 igeblodprovstest
      2 igeförmedlad
      1 igeförmedlade
      1 igelbehandling
      2 igeln
      1 igelns
      1 igemedierad
      2 igemolekyler
    129 igen
      1 igenkännandet
      1 igenkännbar
      2 igenkännbara
      1 igenkännbart
      1 igenkännes
      6 igenkänning
      1 igenkänningsstörningar
      1 igenkänningstecken
     63 igenom
      1 igensatt
      1 igensluten
      2 igetester
     15 igf
      1 igfnivåer
      3 igg
      1 iggantikroppar
      6 iglar
      2 igm
      2 igmantikroppar
      1 ignacio
      6 ignaz
      1 igniarius
      1 ignis
      1 ignorera
      4 ignorerade
      2 ignoreras
      9 ihåg
      1 ihågkommas
      1 ihågkommen
      6 ihålig
      4 ihåliga
      3 ihåligt
     11 ihållande
      1 ihång
      1 ihängande
      3 ihärdiga
      2 ihärdigt
     10 ihjäl
      1 ihjälgasning
      1 ihjälrifven
      2 ihjälriven
    139 ihop
      1 ihopförlänger
      1 ihopklämt
      1 ihopklumpning
      1 ihopkopplade
      1 ihopkurad
      1 ihopläkning
      1 ihoprullad
      1 ihopsydd
      1 ihopväxt
      1 ihopväxta
      1 ihopvirade
      1 ihs
      1 ihsklassifikationen
     51 ii
      1 iia
      1 iialdosteronsystemet
      1 iidiabetiker
     16 iii
      1 i�iii
      1 iiistudier
      1 iireceptorer
      2 iis
      1 iiv
      1 i�iv
      1 ik
      1 ikini
      1 ikke
      1 iklädd
      1 ikon
      1 ikoniska
      9 ikterus
      2 iktus
      2 iktyos
      4 il
      1 ilads
      1 ilägg
      1 iläkemedelskontaminationsymptomen
      7 iländer
      2 iländerna
      1 ilb
      3 ileocekalklaffen
      3 ileostomi
      1 ileostomioperation
      1 ileostomiopererad
      8 ileum
      2 ileus
      1 ilex
      1 iliacakärl
      1 iliotibialbandet
      1 iliotibialbandssyndrom
      1 ilizarovs
      1 ill
     16 illa
      2 illabefinnande
      9 illaluktande
     75 illamående
      1 illamåendedåsighet
      1 illamåenden
      5 illegal
      8 illegala
      4 illegalt
      1 iller
      1 illicium
      1 illinios
      2 illinois
      2 illness
      2 illusion
      1 illusionen
      2 illusioner
      1 illustration
      1 illustrationen
      1 illustrera
      1 illustrerade
      1 illustrerades
      3 illustrerar
      3 illustreras
      1 illvilliga
      1 ilmenium
      2 ilningar
      5 ilo
      1 ilomants
      2 ilos
     10 ilska
      1 ilskan
      2 ilsket
      1 ilskna
      1 iluftvägssekret
      4 im
      1 image
      1 imageskapande
      1 imaginär
      1 imaginära
      2 imaging
      4 imago
      2 imbecilla
      1 imbecillitet
      1 imeretien
      1 imidazolgruppens
      1 imidazolgrupper
      1 imidazolring
      1 imidazopyridinderivat
      1 imigran
      1 imikvimod
      1 imitationer
      1 imitatör
      2 imitatören
      3 imiterar
      1 imiteras
      2 immanuel
      1 immateriellt
      1 immigranter
      2 immitis
      1 immki
      1 immobilisation
      1 immobiliserad
      1 immobiliseras
      1 immortality
      9 immun
     10 immuna
      1 immunadsorberande
      4 immunbrist
      1 immunbrister
      1 immunbristsyndrom
      5 immunbristvirus
      1 immunbristvirusets
      8 immunceller
      1 immuncellerna
      1 immundefekta
      1 immunfixation
      1 immunförsvagad
     59 immunförsvar
     79 immunförsvaret
      6 immunförsvarets
      1 immunförsvarlymfocyterna
      1 immunförsvarret
      1 immunförsvarsaktiveringen
      2 immunförsvarsceller
      1 immunförsvarsreaktion
      1 immunförsvarsrespons
      1 immunglobulin
      1 immunglobulinklass
      1 immunhämmande
      1 immunisera
      6 immunisering
     26 immunitet
      1 immuniteten
      2 immunitetens
      1 immunitetsbildande
      1 immunitetsstatus
      1 immunkomplex
      1 immunkomprometterade
      1 immunmodulerande
      1 immuno
      1 immunoassay
      3 immunodeficiency
      1 immunodeficienta
      1 immunodermatologi
      1 immunofenotypiska
      2 immunofluorescens
      2 immunogena
      1 immunogent
      7 immunoglobulin
      2 immunoglobuliner
      1 immunoglobulinklass
      1 immunoglobulinmolekylerna
      5 immunologi
      1 immunologin
     11 immunologisk
     14 immunologiska
     10 immunologiskt
      1 immunomodulatorer
      1 immunosorbent
      6 immunostimulerande
      1 immunosuppressiv
      1 immunosuppressiva
      1 immunosupprimerade
      1 immunosupressiv
      1 immunosuprimerande
      4 immunoterapi
      2 immunproblem
      2 immunreaktion
      1 immunreaktioner
      2 immunrespons
      2 immunsuppression
      1 immunsuppressiva
      1 immunsuppressivt
      4 immunsupprimerade
      9 immunsvar
      6 immunsvaret
     19 immunsystem
     23 immunsystemet
      7 immunsystemets
      1 immunsystemmodulerande
      7 immunterapi
      1 immuntillstånd
      1 imo
      1 imolekyler
      1 impairment
      2 impedansen
      1 imperativformen
      1 imperatorn
      1 imperfekt
      1 imperial
      1 imperiet
      7 impetigo
     19 implantat
      9 implantaten
      7 implantatet
      1 implantatets
      7 implantation
      1 implantationen
      1 implantatsstorlek
      1 implantatsstorlekarna
      1 implantattekniken
      2 implanterade
      2 implanteras
      1 implantering
      1 implanteringen
      1 implementerandet
      1 implementerar
      1 implementeras
      1 implications
      1 implicerar
      1 implicit
      1 implicita
      1 implikationer
      1 implikationerna
      2 imploderar
      1 implosion
      2 imponerande
      2 import
      1 importaffärer
      1 importerad
      5 importerade
      1 importerades
      5 importeras
      1 importerat
      1 importerats
      1 importör
      2 importören
      1 importörer
     20 impotens
      1 impotenta
      6 impotentia
      1 impregnera
      1 impregnerade
      1 impressionister
      1 impressus
      2 improviserade
     11 impuls
     11 impulsen
      1 impulsens
     22 impulser
      4 impulserna
      1 impulsiv
      3 impulsiva
      8 impulsivitet
      2 impulsiviteten
      1 impulsivt
      3 impulskontroll
     11 impulskontrollstörning
     14 impulskontrollstörningar
      2 impulskontrollstörningarna
      1 impulssignaler
      1 impulsstörningar
      1 impusle
      1 imubakko
    848 in
      1 inackorderingshem
      3 inadekvat
      3 inadekvata
      5 inaktiv
      2 inaktiva
      2 inaktivera
      3 inaktiverade
      2 inaktiverar
      4 inaktiveras
      2 inaktivering
      4 inaktivitet
      1 inaktivitetsatrofi
      2 inaktivt
      3 inälvor
      1 inälvorna
      1 inälvsfasen
      1 inälvsmaskar
      1 inälvsparasit
      1 inälvsparasiter
      1 inandad
      2 inandade
      8 inandas
      1 inandats
     36 inandning
      1 inandningar
      3 inandningen
      1 inandningsgasen
      1 inandningsluft
      4 inandningsluften
      1 inandningsmusklerna
      1 inandningspreparat
      1 inandningsreflex
      2 inandningstryck
      1 inandningstrycket
      2 inari
      1 inarialtare
      1 inärning
     10 inåt
      1 inåtgående
      2 inattentive
      1 inåtuppåt
      1 inåtvänt
      1 inåtväxta
      5 inavel
      1 inavelsproblematik
      1 inbäddad
      2 inbäddade
      1 inbäddat
      3 inbegripa
     14 inbegriper
      1 inbegrips
      3 inbillad
      2 inbillade
      1 inbillar
      1 inbillning
      1 inbillningssjuka
      1 inbindning
      1 inbjöds
      1 inbjudan
      1 inbjudna
      3 inblandad
     27 inblandade
      3 inblandat
      4 inblandning
      3 inblåsningar
      1 inblåsningarmin
      2 inblick
      1 inböjda
      1 inbördes
      1 inbördeskriget
      1 inbringa
      1 inbringat
      1 inbrottslarm
      1 inbrottsskydd
      1 inbunden
      3 inbyggd
      5 inbyggda
      1 inbyggt
      1 inc
      1 incb
      2 incest
      1 inch
      1 inches
      1 incidence
      8 incidens
     11 incidensen
      1 incidensmått
      1 incidenstalen
      3 incidenstalet
      3 incidenter
      1 incidere
      1 incisiverna
      2 incitament
      1 inclusive
      1 inconclusive
      1 inconspicuus
      1 incorporated
      1 incremental
      1 incubus
      1 incurvus
      1 indanderivat
      1 indela
      3 indelad
     27 indelas
      1 indelat
      1 indelkas
     14 indelning
      3 indelningar
      1 indelningarna
      4 indelningen
      1 inden
      1 independent
     10 index
      1 indexera
      1 indexerad
      1 indexerade
      1 indexeringen
      2 india
      2 indiana
      5 indianer
      3 indianerna
      2 indiankulturer
      1 indianskt
      1 indiansstammar
      2 indianstammar
      1 indication
      1 indicators
      3 indicier
      1 indicum
     56 indien
      1 indiens
      1 indier
      1 indifférence
      4 indigo
      1 indigodestillaten
     16 indikation
     15 indikationer
      3 indikationerna
      1 indikationsområden
      1 indikativ
      8 indikator
      3 indikatorer
      1 indikatorerna
      7 indikera
      2 indikerade
      1 indikerande
     23 indikerar
      1 indikeras
      2 indikerat
      1 indir
      1 indira
     18 indirekt
      2 indirekta
     16 indisk
      7 indiska
      2 indiske
      1 indium
     81 individ
      1 individanpassad
     95 individen
     36 individens
      1 individensartens
    191 individer
      6 individerna
      1 individernas
      6 individers
      1 individperson
      1 individplan
      1 individrelaterad
      1 individrik
     10 individs
      1 individtillsynen
      1 individual
      1 individualiseras
      1 individualister
      1 individualistiska
      2 individualitet
      1 individualnivå
     12 individuell
     31 individuella
     28 individuellt
      1 indoeuropeiska
      1 indomalajiska
      1 indometacin
      5 indonesien
      1 indonesisk
      5 indonesiska
      1 indoor
      1 indoprofen
      5 indragen
      2 indraget
      1 indragna
      1 indragning
      1 indränks
      1 indroducerade
      1 induced
      9 inducera
      3 inducerad
      2 inducerade
      1 inducerande
      6 inducerar
      2 induceras
      2 inducerat
      1 inducerbara
      1 induces
      3 induktion
      1 induktionsfas
      2 induktionsfasen
      1 indunstar
      1 indunstas
      3 indunstning
      1 indunstningsresterna
      1 induratum
      1 induseade
      2 induskulturen
     13 industri
      2 industrial
      9 industrialiserade
      1 industrialisering
      2 industrialiseringen
      1 industribagerierna
      1 industribruk
      1 industridesigner
      1 industridesignerna
      1 industridisk
      9 industriell
     10 industriella
     14 industriellt
      2 industrier
      2 industries
      1 industrigrupper
      1 industriguld
      5 industriländer
      4 industriländerna
      1 industrilitteratur
      1 industrilokaler
      1 industrimaten
      1 industrimiljö
     17 industrin
      2 industriöverskott
      2 industrisamhälle
      1 industrisektorn
      1 industriskandalerna
      1 industritomter
      1 industriutsläppen
      1 industrivärlden
      1 industry
      1 ine
      2 ineffektiv
      4 ineffektiva
      1 ineffektivare
      2 ineffektivitet
      3 ineffektivt
      1 inermis
      5 inert
      2 inerta
      1 inertgasens
      1 inevitably
      1 infågande
      1 infälda
      1 infalla
      1 infallande
      5 infaller
      1 infångad
      3 infantil
      1 infärgas
      2 infärgning
     11 infarkt
      3 infarkten
      1 infarkter
      1 infart
      2 infästning
      1 infattar
      1 infattning
      1 infectio
      2 infection
      1 infections
      4 infectious
     19 infektera
     27 infekterad
     82 infekterade
      1 infekterades
      4 infekterande
     16 infekterar
     15 infekteras
     16 infekterat
      9 infekterats
    233 infektion
     95 infektionen
      2 infektionens
    188 infektioner
      4 infektionerna
      1 infektions
      1 infektionsbesvären
      2 infektionsdosen
      1 infektionsduglig
      1 infektionsfallen
      1 infektionsförlopp
      2 infektionsförloppet
      2 infektionsförsvar
      1 infektionsförsvaret
      1 infektionsfrämjande
      2 infektionskänsliga
      3 infektionskänslighet
      2 infektionspsykoser
      2 infektionsrisk
      3 infektionsrisken
     26 infektionssjukdom
     24 infektionssjukdomar
      4 infektionssjukdomen
      1 infektionsskedet
      1 infektionsskyddande
      1 infektionsstället
      1 infektionsstatus
      2 infektionssten
      1 infektionsstenar
      1 infektionssymptom
      1 infektionstakten
      2 infektionstalen
      1 infektionstället
      1 infektionstillfället
      1 infektionstillstånd
      1 infektionsväg
      1 infektionsvägar
      4 infektiös
      5 infektiösa
      5 inferior
      1 inferiora
      1 infertila
     13 infertilitet
      1 infertilitetsproblem
      1 infesta
      1 infestans
      1 infgamma
      1 inficio
      2 infiltrat
      1 infiltration
      1 infiltrationen
      1 infiltrativ
      3 infiltrerar
      1 infinna
      1 infinner
      1 infirmity
      1 inflammatio
    163 inflammation
     35 inflammationen
     24 inflammationer
      1 inflammationerna
      3 inflammationsdämpande
      1 inflammationsdämpning
      1 inflammationsdrivande
      3 inflammationshämmande
      2 inflammationsmarkörer
      1 inflammationsprocess
      1 inflammationsresponssyndrom
      1 inflammationssjukdom
      1 inflammationssjukdomar
      1 inflammationssvar
      2 inflammationssymptom
     21 inflammatorisk
     21 inflammatoriska
      6 inflammatoriskt
      8 inflammerad
     23 inflammerade
      2 inflammeras
      1 inflammerats
      4 inflation
      1 inflationsförsäkring
      1 inflexibla
      2 inflöde
      1 inflödet
      1 influens
     43 influensa
      2 influensaepidemi
      1 influensaepidemier
      1 influensainfektion
      1 influensainfektioner
      9 influensaliknande
     11 influensan
      1 influensapandemi
      2 influensapandemier
      1 influensaprov
      1 influensasäsong
      1 influensasäsongen
      1 influensasmittor
      1 influensasymptom
      3 influensavaccin
      1 influensavaccinering
     24 influensavirus
      1 influensavirusen
      4 influensaviruset
      1 influenser
      2 influenserna
      1 influensor
      1 influensvirus
      1 influenza
     10 influenzae
      1 influenzaemeningit
      1 influerad
      2 influerade
      1 influerades
      1 influerat
     21 inflytande
      1 inflytandet
      5 inflytelserik
      5 inflytelserika
      1 inföll
     76 inför
     14 införa
      7 införande
      1 införandedatum
     14 införandet
      2 införas
      1 införd
      4 införda
     10 införde
     40 infördes
      1 införes
      1 införingshylsa
      1 införlivades
      1 införlivas
      1 införlivats
      1 informatics
    127 information
     17 informationen
      2 informationer
      1 informationsbärande
      1 informationsbehandlande
      1 informationsflödet
      1 informationshjälp
      1 informationskällor
      1 informationskanal
      2 informationskanaler
      1 informationsmaterial
      3 informationsöverföringen
      1 informationssignalerna
      1 informationsspridningen
      1 informationssystem
      1 informationsteknologi
      1 informativa
      2 informell
      4 informella
      1 informellt
      7 informera
      2 informerad
      1 informerar
      1 informeras
      2 informerat
      6 införs
      4 införsel
      1 införseln
      1 införseltillstånd
      2 införskaffa
      4 infört
      8 införts
      1 infraljud
      1 infraröda
      2 infrarött
      2 infrastruktur
      1 infrastrukturen
      2 infrusen
      1 infrysning
      1 infryst
      1 infundibulum
      6 infusion
      1 infusioner
      1 infusionssalt
      1 infusionsvätska
    151 inga
     24 ingå
     13 ingående
      3 ingång
      6 ingången
      1 ingångsporten
      1 ingångssäkringarelmätare
      1 ingångsspalt
      1 ingångsställe
    152 ingår
      1 ingås
      2 ingått
      2 inge
      1 ingeborg
      1 ingelman
      1 ingemansson
      1 ingemar
    238 ingen
      2 ingendera
      1 ingenjör
      1 ingenjören
      1 ingenjörskonsten
      7 ingenting
      1 ingestion
    108 inget
      1 ingetdera
      1 ingett
      3 inghe
     18 ingick
      1 ingivelse
      1 ingivelser
      1 inglasade
      1 ingram
      9 ingrediens
      1 ingrediensen
      8 ingredienser
      3 ingredienserna
      1 ingredient
     93 ingrepp
      4 ingreppen
     25 ingreppet
      1 ingreppetref
      4 ingripa
      6 ingripande
      1 ingriper
      1 ingrupperas
      1 ingvar
      1 inh
      2 inhägnad
      1 inhägnade
      1 inhägnat
      2 inhalation
      1 inhalationen
      2 inhalationsanestesi
      2 inhalationsform
      1 inhalationsinduktion
      1 inhalationsläkemedlet
      3 inhalationsmedel
      3 inhalationsnarkos
      4 inhalationssteroid
      5 inhalationssteroider
      1 inhalationssteroidlångverkande
      4 inhalator
      1 inhalatorer
      2 inhalatorn
      2 inhalera
      1 inhalerande
      3 inhaleras
      1 inhalering
      3 inhämta
      1 inhämtar
      3 inhämtas
      1 inhandla
      1 inhandlades
      3 inhemsk
      2 inhemska
      5 inhibera
      1 inhiberade
      1 inhiberande
      3 inhiberar
      1 inhibering
      1 inhibition
      1 inhibitionsbeslutet
      2 inhibitor
      1 inhibitorer
      3 inhibitoriska
      1 inhumant
      1 inhyrd
      1 ini
      1 iniativtagarna
      5 inifrån
      3 initial
      6 initiala
      1 initialern
      2 initialskedet
     15 initialt
      1 initiationsrit
      7 initiativ
      2 initiative
      1 initiativet
      1 initiativförmåga
      1 initiativförmågan
      3 initiativlöshet
      2 initiera
      1 initierade
      2 initierar
      4 initieras
      1 initierat
      1 injaga
     32 injektion
      2 injektionen
     15 injektioner
      1 injektioninfusion
      1 injektionsbehandling
      2 injektionsform
      1 injektionskanyler
      1 injektionsmissbruk
      1 injektionsnål
      1 injektionsområdet
      1 injektionsredskap
      2 injektionsspruta
      5 injektionsstället
      1 injektionsvätska
      1 injektionsvätskor
      5 injektionsverktyg
      1 injektorer
      6 injicera
      2 injicerade
      1 injicerades
      3 injicerande
      6 injicerar
     13 injiceras
      2 injicerat
      1 injicerats
      1 injicerbara
      1 injicering
      1 inka
      1 inkafolket
      1 inkaindianerna
      1 inkallande
      1 inkallelsebränningar
      1 inkapabel
      1 inkapslad
      1 inkapslade
      2 inkapslat
      1 inkarnerad
      1 inkl
      1 inklämning
      1 inklämt
     12 inkludera
      1 inkluderade
      5 inkluderande
     81 inkluderar
     11 inkluderas
      8 inkluderat
      1 inkluderats
      1 inkludering
      2 inklusions
      2 inklusionskriterierna
      3 inklusionskroppsmyosit
     85 inklusive
      1 inkoherens
      1 inkoherent
      8 inkommande
      1 inkommit
      1 inkomna
      1 inkompetens
      3 inkomplett
      1 inkomst
      3 inkomster
      1 inkomstkällorna
      1 inkomstskillnader
      2 inkonsekventa
     16 inkontinens
      1 inkontinenshjälpmedel
      1 inkontinensproblemen
      5 inkontinensskydd
      1 inkontinensvård
      1 inköp
      1 inköpare
      1 inkopplad
      2 inkopplade
      1 inkopplades
      1 inköpta
      1 inköpte
      1 inköptes
      1 inkorporation
      2 inkorporera
      1 inkorporerad
      1 inkorporerade
      1 inkorrekta
      2 inkörsport
      1 inkräktande
      1 inkräktare
      1 inkringliggande
      1 inkubation
      1 inkubationsfas
      1 inkubationsperioden
     15 inkubationstid
     32 inkubationstiden
      1 inkubator
      1 inkuberar
      1 inkuberingen
      2 inkvisitionen
      3 inkvisitionens
      1 inkvisitor
      1 inkvisitorerna
      4 inlagd
      7 inlagda
      1 inlägg
     10 inläggning
      1 inläggssula
      1 inlagras
      3 inlagring
      1 inlagringen
      2 inlämnades
      2 inland
      2 inlandet
      2 inlandstaipan
      8 inlandstaipanen
      2 inlärd
      4 inlärda
     17 inlärning
      2 inlärningen
      1 inlärningsfaktorer
      2 inlärningsförmåga
      1 inlärningsmekanismen
      1 inlärningsperiod
      1 inlärningsprocesser
      1 inlärningspsykologi
      1 inlärningssituation
      7 inlärningssvårigheter
      1 inlärningsteoretisk
      1 inlärningsteoretiska
      2 inlärningsteori
      6 inleda
      9 inledande
      4 inledas
      2 inledde
      5 inleddes
      1 inleder
      3 inledning
      2 inledningen
      1 inledningsfasen
     13 inledningsvis
     19 inleds
      1 inlemma
      1 inlemmade
      1 inlemmas
      1 inlemmats
      1 inlett
      1 inletts
      2 inlevelse
      1 inlevelseförmågan
      1 inlösen
      1 inmärkt
      1 inmottagningar
      1 inmundigandet
    313 innan
      2 innandöme
     13 innanför
      1 innanpåliggande
      3 innat
      1 innata
     48 inne
     19 innebar
    604 innebär
     40 innebära
      2 innebärande
      1 innebärt
      4 inneboende
      8 innebörd
      4 innebörden
      1 innebörder
      9 inneburit
     12 innefatta
      2 innefattade
      1 innefattades
      3 innefattande
    102 innefattar
      6 innefattas
      1 innefattat
      1 innefattats
      1 innefinner
      1 inneftattar
      9 inneha
     40 innehåll
     40 innehålla
     39 innehållande
      1 innehållandes
    311 innehåller
     15 innehållet
      1 innehållets
      4 innehållit
      2 innehållsämnen
      1 innehållsfilter
      1 innehållsförteckningar
      2 innehållsförteckningen
      1 innehållslös
      1 innehållsstörning
      1 innehållsstörningar
      8 innehar
      2 innehas
      7 innehav
      1 innehavaren
     18 innehöll
      5 inneliggande
      1 inner
      2 innerdiameter
      1 innerkant
      7 innerörat
      1 inneröronens
      2 innerst
      3 innersta
      2 innervägg
      1 innerväggar
      1 innervation
      1 innervävnader
      1 innerverande
      3 innerverar
      2 innerveras
      1 innerveringen
      2 innesluta
      4 innesluten
      4 innesluter
      1 inneslutet
      4 inneslutna
      1 innevarande
      3 innovation
      1 innovationer
      1 innovativ
      1 innovatoinerna
      1 innsbruck
      1 inofficiell
      2 inofficiella
      1 inokulation
      1 inokuleras
   1081 inom
     17 inomhus
      1 inomhusblommor
      1 inomhuscentrum
      1 inomhusluft
      1 inopererad
      1 inordnas
      1 inosilikater
      1 inositol
      1 inpå
      1 inpackning
      1 inpackningar
      1 inpassa
      1 inpassning
      1 inplantera
      1 inplanterade
      1 inplanteras
      1 inplanterat
      1 inpräntade
      1 input
      2 inputs
      1 inquiry
      2 inräknade
      2 inräknar
      2 inräknas
      2 inräknat
      2 inrapporterade
      5 inrätta
      1 inrättad
      1 inrättade
     11 inrättades
      2 inrättande
      1 inrättas
      1 inrättats
      2 inrättning
      2 inrättningar
    124 inre
      1 inreddes
      1 inredning
      1 inredningstextilier
      1 inrepp
      1 inrikes
      1 inrikesflygplanet
      1 inrikta
     11 inriktad
      7 inriktade
      3 inriktar
      7 inriktas
      2 inriktat
      1 inriktats
     24 inriktning
      3 inriktningar
      2 inriktningarna
      4 inriktningen
      1 inrymde
      1 inrymmer
      1 inrymt
     11 insåg
      1 insamla
      2 insamlade
      2 insamlas
      1 insamlats
      1 insamling
      1 insamlingar
      1 insamlingsexpeditioner
      1 insamlingsmetod
      1 insändare
      1 insändes
      1 insane
      1 insanity
      8 insats
      2 insatsen
     47 insatser
     10 insatserna
      1 insatsstyrkan
      1 insatstiden
      1 insatstider
      1 insatstiderna
      1 insatsvärde
      3 insatt
      5 insättande
      1 insättandet
      6 insättning
      5 insätts
      1 insatyrkan
      1 inscribe
      7 inse
      5 insekt
      3 insekten
     35 insekter
      1 insekterdet
      6 insekterna
      1 insektförutom
      1 insektgift
      1 insekticid
      2 insektsangrepp
      1 insektsätare
      2 insektsbekämpning
      5 insektsbett
      1 insektsbiologin
      1 insektsburen
      3 insektsgift
      2 insektsgifter
      1 insektsgruppen
      5 insektsmedel
      1 insektsmedlet
      2 insektsordningen
      1 insektspollinerade
      1 insektsproblem
      1 inseminare
     16 insemination
      3 inseminationen
      1 inseminationer
      1 inseminatus
      1 inseminera
      2 inseminering
      1 insensitivitet
      3 inser
      2 insett
     15 insida
     27 insidan
      1 insidor
      5 insignalen
      2 insignier
     10 insikt
      2 insikten
      6 insikter
      3 insipidus
      1 insituet
      1 insjöar
      8 insjukna
     27 insjuknade
     16 insjuknande
      1 insjuknandefrekvensen
      2 insjuknanden
     16 insjuknandet
     28 insjuknar
      7 insjuknat
      1 insjunkna
      1 inskjutna
      1 inskjuts
      4 inskränker
      2 inskränkning
      1 inskränkningar
      1 inskränkta
      1 inskränktes
      1 inskriven
     29 inslag
      2 inslagen
      1 inslaget
      1 insmord
      1 insmörjningar
      1 insmort
      1 insnitt
      1 insnittet
      6 insomnande
      7 insomni
      1 insomnia
      1 insöndrande
      1 insöndrar
      4 insöndras
      1 insöndring
      2 insöndringen
      3 inspektera
      1 inspekteras
      4 inspektion
      5 inspektionen
      2 inspektioner
      1 inspelade
      1 inspelning
      1 inspelningen
      1 inspelningselektrod
      4 inspiration
      1 inspirationen
      1 inspirationskälla
      2 inspirerad
      2 inspirerade
      1 inspirerades
      1 inspireras
      2 inspirerat
      3 inspirerats
      1 insprirerad
      1 insprutat
      5 instabil
      5 instabila
      3 instabilitet
      1 instabilt
      1 inställd
      1 inställda
      3 inställer
      1 installera
      3 installerad
      1 installerade
      2 installerades
      2 installeras
      1 installerat
      3 installerats
      8 inställning
      3 inställningar
      1 inställningen
      1 inställsamhet
      1 inställt
      1 instängd
      1 instängda
      3 instans
      5 instanser
      1 instickningen
      2 instiftade
      3 instiftades
      5 instinkter
      1 instinkthandlingar
     13 institut
     18 institute
      1 instituten
     26 institutet
      2 institutets
      9 institution
      1 institutionalisera
      1 institutionaliserades
      1 institutionaliserar
      1 institutionella
      7 institutionen
      9 institutioner
      3 institutionerna
      1 institutioners
      1 institutionsvård
      1 instituto
      1 instruera
      1 instruerade
      1 instruerar
      1 instrueras
      9 instruktioner
      4 instruktionerna
      1 instruktionstekniken
      1 instruktörer
    121 instrument
      1 instrumentala
      1 instrumentalsträngar
      1 instrumentalt
      2 instrumentell
      2 instrumentella
     13 instrumenten
      1 instrumenter
     31 instrumentet
      6 instrumentets
      2 instrumentmakaren
      1 instrumentpaneler
     11 insufficiens
      1 insugen
      5 insula
      1 insulatard
     73 insulin
      1 insulinbehandlade
      1 insulinbehov
      1 insulinberoende
      2 insulinbrist
      2 insulinbristen
      1 insulinceller
      1 insulinchocker
      1 insulinderivat
      1 insulindosering
      1 insuliner
     14 insulinet
      2 insulininjektion
      3 insulininjektioner
      1 insulinkänning
      2 insulinkänningar
      2 insulinkänslighet
      2 insulinkoma
      1 insulinkomabehandling
      1 insulinkrävande
      1 insulinlike
      1 insulinliknande
      2 insulinmolekylen
      4 insulinnivåer
      1 insulinnivån
      1 insulinpåslaget
      2 insulinproducerande
      1 insulinproduktionen
      2 insulinpump
      1 insulinpumpar
      4 insulinpumpen
      1 insulinreceptorer
      6 insulinresistens
      1 insulinsorter
      1 insulintillförsel
      1 insult
      1 insuman
      1 insydda
      2 insyn
      8 inta
     66 intag
      4 intåg
      4 intagande
      2 intagandet
      2 intagas
      2 intagen
      4 intages
     17 intaget
      4 intagit
      9 intagits
      3 intagna
      8 intakt
      5 intakta
      3 intäkter
      1 intäkterna
      1 intala
     14 intar
     22 intas
   3726 inte
      1 integralt
      1 integras
      3 integrated
      2 integration
      2 integrera
      3 integrerad
      3 integrerade
      1 integrerades
      1 integrerande
      6 integrerar
      2 integreras
      2 integrerat
      1 integreringsprocessesen
      4 integritet
      1 integriteten
      1 intellego
      2 intellekt
      2 intellektet
      1 intellektualism
      6 intellektuell
     11 intellektuella
      4 intellektuellt
      3 intelligence
     48 intelligens
      3 intelligensbegreppet
      1 intelligensbrist
      9 intelligensen
      1 intelligensens
      2 intelligenser
      1 intelligensfaktor
      1 intelligensforskning
      6 intelligenskvot
      1 intelligenskvoten
      1 intelligensmätning
      1 intelligensmätningen
      3 intelligensnivå
      1 intelligensprofil
      1 intelligensprofiler
      1 intelligensteori
      4 intelligenstest
      2 intelligenstesten
      2 intelligenstester
      1 intelligenstestet
      1 intelligent
      3 intelligenta
      1 intelligenzquotient
      1 intensifieras
      1 intensifierat
      1 intensifiering
     18 intensitet
     33 intensiv
     14 intensiva
      3 intensivare
      1 intensive
     11 intensivt
     14 intensivvård
      3 intensivvården
      3 intensivvårdsavdelning
      3 intensivvårdsavdelningar
      1 intensivvårdsavdelningreceptfri
      1 intensivvårdsenhet
      1 intensivvårdsinsats
      1 intensivvårdsläkare
      1 intensivvårdssjuksköterska
      1 intention
      1 intentionalitet
      2 intentioner
      1 interacting
      3 interaction
      7 interagera
      5 interagerar
     12 interaktion
      5 interaktionen
     10 interaktioner
      1 interaktionerna
      1 interaktionsfärdigheter
      1 interaktionsrisk
      1 interarytenoidmuskel
      3 intercostales
      1 intercostalmuskulatur
      1 interdentalborste
      1 interdiciplinärt
      1 interdigestivfasen
      1 interdigital
      1 interdisciplinära
      3 interferon
      5 interferoner
      2 interimanalys
      1 interimanalyser
      1 interindividuella
      1 interkontinentala
      1 interleukin
      1 interleukiner
      1 intermedia
      1 intermediär
      1 intermediärer
      1 intermediat
      2 intermittens
      9 intermittent
      1 intermolekylära
      4 intern
     11 interna
      1 internal
      1 internaliseras
     22 international
      1 internationale
     18 internationell
     58 internationella
     47 internationellt
      1 interner
     22 internet
      1 internetanvändning
      1 internetbaserat
      1 internetbehandling
      2 internetberoende
      1 internetenkät
      1 internetforum
      1 internetforumet
      1 internethistorik
      1 internets
      1 internetsidan
      1 internetsidor
      1 internetspel
      2 internetterapi
      1 internettrafik
      2 interneuron
      2 interni
      1 internkontroll
      2 internmedicin
      1 internmedicinare
      1 internordiska
      2 internt
      1 internus
      1 internutredning
      1 interoception
      2 interpersonell
      1 interpunktion
      1 interstellära
      1 interstitialcell
      1 interstitialvätska
     17 interstitiell
      1 interstitiella
      1 interstitiellt
      1 intersubjektivitet
     14 intervall
      1 intervallbehandling
      2 intervaller
      7 intervallet
      1 intervallträning
      1 intervenera
      1 intervenerade
      1 intervension
     10 intervention
      1 interventionen
      6 interventioner
      1 intervertebraldiskarna
      1 interview
      2 interviewrevised
      2 intervju
      1 intervjua
      2 intervjuades
      1 intervjuar
      1 intervjubaserad
      1 intestinala
      1 intestinalmetaplasi
      3 intestinum
      2 intet
      1 intetsägande
      1 inti
     21 intill
     15 intilliggande
      3 intim
      3 intima
      1 intimrakning
      5 intimt
      1 intöcknande
      2 intog
      4 intolerans
      1 intoleranser
      1 intoxikation
      2 intoxikationer
      2 intra
      1 intraabdominellt
      1 intraartikulär
      1 intracellulär
      8 intracellulära
      6 intracellulärt
      4 intracerebral
      1 intracervical
      3 inträdde
      4 inträde
     18 inträder
      1 inträdet
      1 intraepiteliala
     31 inträffa
     28 inträffade
     56 inträffar
     17 inträffat
      1 intrahepatiska
      2 intrakavitär
      2 intrakraniell
      4 intrakraniella
      7 intrakraniellt
      2 intramuskulär
      1 intramuskulära
      4 intramuskulärt
      1 intrång
      1 inträngade
      1 inträngandet
      1 inträngt
      1 inträning
      2 intraokulära
      1 intraokulärt
      1 intraperitoneal
      1 intrapersonell
      1 intratekal
      1 intratekalt
      1 intrathekal
      1 intratorakala
      5 inträtt
      4 intrauterin
      1 intrauterina
      1 intravaginala
      2 intravasal
     21 intravenös
      8 intravenösa
     29 intravenöst
      1 intravenöstvårdpersonal
     14 intressant
      3 intressanta
     31 intresse
      3 intressebevakningsfullmakt
      1 intresseförening
      3 intresseföreningar
      4 intressen
      3 intressenter
      1 intresseområden
      1 intresseorganisation
      2 intressera
      9 intresserad
      4 intresserade
      2 intresserar
     19 intresset
      1 intriger
      1 intrikata
      2 intrinsic
      1 intrinsikalt
      2 intrinsiska
     19 introducerade
     26 introducerades
      1 introducerar
      2 introduceras
      5 introducerats
      6 introduktion
      2 introduktionen
      1 introduktionskurs
      1 introlåt
      1 intrusiva
     11 intryck
      3 intrycken
      5 intrycket
      3 intryckt
      8 intubation
      2 intubera
      1 intuberad
      1 intuberas
      2 intubering
      1 intuition
      1 intuitiv
      1 intuitiva
      2 intussusception
      1 intyg
      2 inuiterna
      2 inuiternas
      1 inulin
     59 inuti
      7 invadera
      6 invaderar
      3 invaderas
      2 invagination
      2 invalider
      2 invalidiserade
      2 invalidiserande
      3 invaliditet
      1 invånarantalet
     17 invånare
      5 invånarna
      3 invanda
      1 invänder
      1 invändig
      7 invändigt
      1 invändningar
      1 invandrade
      3 invandrare
      1 invandrargrupper
      1 invandring
      1 invänt
      2 invänta
     11 invärtes
      3 invärtesmedicin
      3 invärtesmedicinska
      6 invasion
      1 invasionen
      1 invasionshärar
     15 invasiv
     12 invasiva
      2 invasivt
      1 inväxta
      2 invecklade
      2 inventering
      1 inventeringar
      1 inventory
      2 inverka
      1 inverkade
     51 inverkan
     10 inverkar
      1 inversion
      2 inverterade
      1 inverterat
      5 investera
      1 investerar
      1 investerare
      1 investerat
      5 investering
      4 investeringar
      1 investeringarna
      1 investeringen
      1 investeringsguld
      4 invid
      2 inviga
      1 invigd
      2 invigdes
      1 invivider
      1 involutus
      2 involvera
     13 involverade
     23 involverar
      3 involverat
      1 inwriteto
      1 inympas
      1 iode
      1 iodes
      1 iodine
      3 iögonfallande
      1 iohexol
      2 iom
      1 ion
      1 ionisation
      1 ionization
      1 ionizing
      2 iop
      1 iowa
      1 ipa
      1 ipbaserad
      1 ipccs
      1 iphone
      2 ipratropium
      4 ips
      4 ipseo
      1 ipsilaterala
      1 ipsilateralt
      1 ipt
     35 iq
      1 iqföreningar
      1 iqnivån
      1 iqpoäng
      5 iqtest
      4 iqtester
      2 iqvärde
      1 iqwig
      1 ir
      3 irak
      1 irakkriget
     11 iran
      1 iranska
      1 ireceptorer
      1 irgasan
      1 iridektomi
      1 iridium
      1 iridologin
     21 iris
      1 irisdiagnostik
      1 irisdiagnostiken
      1 irisdiagnostikens
      3 irisen
      1 irish
      1 irisheterokromi
      2 irisin
      1 irisoch
      1 iristopografi
      1 irisvävnaden
     10 irit
      2 iriter
     22 irland
      1 irlands
      1 irländsk
      1 irländska
      1 iron
      1 ironbinding
      1 ironiskt
      1 irrar
      3 irrationell
      2 irrationella
      2 irrationellt
      1 irrelevant
      4 irrelevanta
      1 irreparabel
      1 irreversibel
      1 irreversibelt
      1 irreversibla
      1 irrigation
      5 irritabel
      4 irritabilitet
      1 irritans
      1 irritanter
     17 irritation
      1 irritationer
      1 irritationlokala
      1 irritera
      2 irriterad
      1 irriterade
     14 irriterande
      6 irriterar
      3 irriteras
      1 irrlära
      1 irstrålning
      3 irukandji
      1 irukandjimaneten
      1 irving
     16 is
      1 isaa
      2 isaac
      2 isabella
      2 isadora
      1 isak
      1 isande
      4 isär
      1 isättika
      1 isbad
      1 isberg
      1 isbjörn
      3 isbn
      1 iscensättningar
     10 ischemi
      1 ischemin
      6 ischemisk
      1 ischemiska
      5 ischias
      2 ischiasnerven
      2 ischiasnervens
      1 ischnocera
      2 isen
      1 isens
      1 isfolket
      1 isformationer
      1 ishacka
      1 ishockeyspelare
      1 isigt
      1 isigtsnöigt
      1 ising
      1 iskall
      1 iskariot
      2 iskristaller
      1 isl
      1 isla
      5 islam
      1 islamiska
      1 islamistiskpalestinska
      2 islams
      4 island
      2 isländska
      1 isländskans
      3 ismannen
      2 isningar
      3 iso
      1 isocyanater
      1 isoelektriska
      2 isoenzymer
      3 isofluran
      1 isogami
      3 isoinokosteron
      1 isolat
      1 isolation
      1 isolationsmaterial
     15 isolera
      4 isolerad
     11 isolerade
      6 isolerades
      2 isolerande
      8 isolerar
      7 isoleras
      8 isolerat
      2 isolerats
     31 isolering
      1 isoleringens
      1 isoleringsåtgärder
      1 isoleringseffekt
      1 isoleringsmaterial
      4 isomer
      1 isomera
      1 isomeren
      1 isomerer
      1 isomererna
      1 isomerpar
      1 isomorft
      1 isonandra
     10 isoniazid
      1 isoosmolär
      3 isopati
      2 isopatin
      2 isopropanol
      1 isopropylalkohol
      1 isopropylbensen
      1 isopropylmetakresol
      1 isopropylmetylfenol
      1 isopropylmetylfluorfosfonat
      1 isostandard
      6 isotop
     13 isotopen
      5 isotoper
      1 isotophalterna
      1 isotopmärkta
      1 isotopundersökning
      1 isoxapenicilliner
      1 isoxapenicillinerna
      1 isoxazolylpenicilliner
      1 ispåse
      7 israel
      1 israelisk
      4 israeliska
      1 israeliter
      1 israeliterna
      2 israels
      2 issykkul
    220 istället
      1 ister
      2 isthmus
      2 istiden
      3 it
      2 itaa
      1 itaas
     40 italien
      1 italienborg
      2 italiensk
     10 italienska
      2 italienskans
      2 italienske
      1 italienskt
      1 itinfrastrukturs
      1 itis
      4 itp
      1 itrakonazol
      3 its
      2 itstress
      6 itu
      3 iucn
      1 iucns
      3 iupac
      3 iupacnamn
      1 iutrymme
     17 iv
      1 iva
      7 iväg
      2 ivan
      1 ivd
      2 ivermectin
      2 ivf
      3 ivo
      2 ivory
      1 ivrigt
      3 ivy
      1 ivydermatit
      2 ivymetoden
      1 iwakami
      1 i[williamsburg
      7 ix
      1 ixodes
      1 [ixodes
      1 iyengar
      1 iyengaryoga
     13 j
      9 ja
      1 jack
      2 jackins
      1 jackor
      7 jackson
      2 jacksons
      2 jacob
      3 jacobs
      1 jacq
      4 jacques
      2 jadad
      1 jadadbechara
      2 jadadskalan
      2 jade
     16 jag
      3 jaga
      3 jagade
      5 jagar
      2 jägar
      6 jägare
      1 jägaren
      1 jägaresamlare
      1 jägarfolk
      1 jägarliv
      3 jägarna
      2 jagas
      1 jagdrifterna
      1 jagellonica
     20 jaget
      1 jagetsjälen
      1 jagfunktion
      1 jagfunktionen
      6 jagfunktioner
      2 jagfunktionerna
      1 jagkänsla
      4 jagpsykologin
      1 jagpsykologiska
      1 jagstyrd
      9 jakob
     11 jakt
      1 jäkt
      1 jakten
      1 jaktlagar
      1 jaktlyckan
      1 jaktstuga
      1 jaktvapen
      1 jalappa
      1 jama
      1 jamahl
      1 jämbördigt
     18 james
     38 jämför
     15 jämföra
      3 jämförande
     17 jämföras
      4 jämförbar
      3 jämförbara
      2 jämförbart
      3 jämförde
      4 jämfördes
      1 jämförels
     21 jämförelse
      1 jämförelsegrupper
      1 jämförelsemått
      2 jämförelsen
      5 jämförelser
      4 jämförelsevis
      6 jämförs
     90 jämfört
      1 jämförts
      1 jämlikhetsaspekter
     14 jämn
     12 jämna
      1 jämnar
      1 jämnare
      5 jämnåriga
      2 jämnas
      1 jämnstora
      6 jämnt
      1 jämnvarma
      1 jämställde
      4 jämställdhet
      1 jämställdheten
      1 jämställdhetsaspekter
      1 jämställer
      1 jämställs
      3 jämställt
      1 jämställts
      2 jämte
      2 jämtland
      1 jämtlands
      9 jämvikt
      2 jämvikten
      1 jämviktsförhållande
      1 jämviktsnivå
      7 jan
      1 janakananda
      8 janet
      1 janez
      3 jani
      1 janis
      1 janne
      6 janov
      3 janovs
      1 jansdotter
     33 januari
      1 jap
     45 japan
      1 japanen
      2 japaner
      2 japans
      8 japansk
     24 japanska
      1 japanskan
      1 japanske
      2 japanskt
      3 japonicus
      1 jared
      1 jari
     36 järn
      1 järna
      1 järnaffärer
      1 järnålder
      5 järnåldern
      4 järnatomen
      1 järnatomens
      1 järnbärande
      1 järnberikade
      1 järnbeslag
      7 järnbrist
      1 järnbromid
      3 järndepåer
      1 järndepåerna
      3 järnet
      1 järniiiklorid
      1 järniijoner
      1 järn[ii]oxygenoxidoreduktas
      1 järnindustri
      1 järninnehållande
      2 järnjon
      1 järnkälla
      2 järnklorid
      1 järnklump
      1 järnlunga
      1 järnlungan
      1 järnmättnad
      1 järnmetabolismen
      2 järnnivåer
      7 järnöverskott
      1 järnskenor
      1 järnspisens
      1 järnstatus
      1 järnsulfat
      1 järntillskott
      1 järntransportproteinet
      1 järntribromid
      1 järnupptag
      1 järnupptaget
      3 järnväg
      1 järnvägarna
      5 järnvägen
      1 järnvägsbygge
      1 järnvägsetablering
      4 järnvägskorsning
      1 järnvägskorsningar
      1 järnvägsövergångarna
      1 järnvägsspår
      1 järnvägsstation
      1 järnvägstrafik
      1 järnvägsvagnar
      1 järnvärcktyg
      1 jaröster
      1 järv
      1 järvsö
      1 jäsbar
      1 jäser
      5 jäsning
      1 jäsningen
      1 jäsningsprocess
      2 jäsningsteknologi
      4 jaspers
      1 jäst
      1 jäste
      2 jästen
      1 jästkulturer
      1 jästliknade
      6 jastreboff
      3 jästsvamp
      2 jästsvampar
      1 jästsvamparna
      2 jästsvampen
      1 jätte
      1 jättebjörnloka
      3 jättebjörnlokan
      1 jättebläckfisken
      2 jätteceller
      4 jättecellstumör
      5 jätteloka
      2 jättelokan
      1 jättelokor
      1 jättelokorna
      1 jättenysrot
      1 jätteproppen
      1 jättestor
      1 jättestorlek
      1 jätteticka
      1 jättetickan
      1 jättetonsilloliter
      3 jättevaran
      3 jättevaranen
      1 jättevarg
      4 jätteväxt
      1 jäv
      1 java
      2 javel
      1 javelle
      1 jävig
      1 jay
      1 jaye
      1 jaynes
      1 jazz
      1 jb
      1 jbs
      2 je
      6 jean
      2 jeanbaptiste
      1 jeancharlesmarcantoine
      1 jeanfran�ois
      1 jeanmarc
      1 jeans
      1 jeff
      4 jehovas
      1 jejunostomi
      4 jejunum
      1 jekyll
      1 [jenes]
      8 jenner
      1 jennifer
      1 jens
      2 jensen
      1 jepsonii
      1 jeremias
      1 jerker
      1 jeronimo
      1 jerrys
      5 jersey
      2 jerusalem
      1 jerusalemsyndromet
      1 jerzy
      1 jesaja
      3 jesu
      1 jesuiten
     11 jesus
      1 jesusbarnet
      1 jetflygplan
     11 jetlag
      1 jetpacks
      1 jetplan
      1 jf
      3 jfr
      1 jihad
      1 jim
      2 jimi
      1 jindynastin
      1 jiroveci
      1 jivamuktiyoga
      1 jivan
      1 jivanmukta
      1 jivatma
      1 jk
      1 jkg
      3 jmf
      2 jmfr
      1 jnanayoga
      1 joachim
      1 joan
      6 jobb
      7 jobba
      3 jobbade
      9 jobbar
      1 jobbat
      1 jobben
     12 jobbet
      1 jobbiga
      2 jobbigt
     43 jod
      2 jodatomer
      1 jodbasedows
      1 jodberikat
      7 jodbrist
      1 jodbristsyndrom
      1 joderingsprogram
      1 jodfenol
      2 jodföreningar
      2 jodförgiftning
      1 jodhaltigt
      3 jodid
      1 jodiden
      1 jodidjoner
      1 jodidlösningar
      2 jodie
      3 jodkalium
      3 jodkälla
      1 jodkällorna
      2 jodlösning
      6 jodmetan
      6 jodoform
      1 jodoformens
      1 jodoformtestet
      2 jodsyrat
      1 jodtillskott
      1 jodtyrosindejodinas
      1 joe
      1 joel
      9 johan
      4 johann
      1 johanna
      4 johannes
      1 johannesberg
      2 johannisson
     13 johansson
     37 john
      1 johnny
      2 johns
      1 johnson
      1 johnsons
      2 joint
      1 jointar
      1 jois
      1 jojoba
      1 jok
      1 jolt
      4 jon
      1 jón
      3 jonas
      3 jonathan
      1 jonbalans
      1 jonbytare
      1 jonbyte
      1 jonen
     20 joner
      5 jonerna
      1 jonernas
      1 joners
      2 jonfälla
      3 jonförening
      1 jonglera
      1 jongradienter
      3 joniserade
     24 joniserande
      1 joniserar
      1 joniseras
      5 jonisering
      1 joniseringssystem
      1 jonium
      2 jonkanal
     14 jonkanaler
      3 jönköping
      1 jönköpings
      1 jonlösning
      1 jonotropa
      1 jonpumpar
      1 jonpumparna
      1 jöns
      3 jonsson
      1 jonströmmar
      1 jonvikt
     28 jord
      2 jordabalken
      1 jordanien
      2 jordar
      1 jordarter
      3 jordartsmetaller
      1 jordartsmetallerna
      1 jordbävning
      3 jordbävningar
      1 jordbävningen
      4 jordbruk
      1 jordbrukare
      5 jordbruket
      2 jordbrukets
      2 jordbruksmark
      1 jordbruksorganisation
      2 jordbruksprodukter
      1 jordbrukssamhället
      1 jordbrukssamhällets
      2 jordbruksutveckling
      1 jordbruksutvecklingsfonden
      1 jordbruksverk
      3 jordbruksverket
      1 jordbruksverks
      4 jorddragning
      2 jorddragningen
      1 jordegumma
      1 jordegumman
      1 jordegummorna
      2 jordekorrar
      1 jordelektrod
      1 jordeliv
      1 jordelivet
      1 jordemoder
      4 jordemodern
      2 jordemödrarna
      7 jordemor
      1 jordemorbarnmorska
      1 jordemorskrået
     33 jorden
     17 jordens
      3 jordfast
      1 jordfilter
      1 jordgubben
      1 jordgubbsplantorna
      1 jordgumma
      2 jordgumman
      1 jordhögar
      1 jordisk
      1 jordiska
      1 jordmor
      1 jordnöts
      6 jordnötsallergi
      1 jordnötsallergiker
     13 jordnötter
      1 jordreva
      4 jordrök
      1 jordröken
      1 jordröksväxter
      1 jordskiktet
      5 jordskorpan
      6 jordstam
      2 jordstammar
      3 jordstammen
      1 jordstammens
      1 jordtyper
      2 jordytan
      2 jörgen
      2 josé
      2 josef
      2 josefsson
     12 joseph
      1 josephine
      1 jössel
      3 joule
      1 jourmottagningar
     22 journal
      2 journalen
      4 journaler
      1 journalföring
      1 journalist
      2 journalisten
      1 journalister
      2 journalsystem
      1 joyce
      1 j�rgen
     74 ju
      1 juan
      1 jubileumssanatorier
      1 juda
     13 judar
     10 judarna
      1 judarnas
      2 judas
      1 judeförföljelsen
      1 judeförföljelser
      1 judehat
      1 judehatet
      2 judendomens
      4 judiska
      1 judith
      2 judo
      2 juice
      1 julbadet
      1 julep
      3 jules
      1 julesÉmile
      1 julhelgen
     27 juli
      1 julia
      2 julian
      1 juliaugusti
      1 juli�augusti
      4 julius
      1 julpyntning
      1 julros
      1 julrosen
      1 julrosor
      2 julrosorna
      1 julrossläktet
      2 julstädning
      1 junctions
      1 jünger
      2 jungfrufödsel
      2 jungfrun
     30 juni
      2 juniaugusti
      4 junijuli
      1 junin
      1 juniperus
      1 junktursignal
      1 jurabergen
      1 jurgens
      4 juridik
      4 juridisk
      3 juridiska
     14 juridiskt
      2 jurisdiktion
      1 jurisdiktioner
      2 jurist
      1 juryn
      1 jusjtjenko
      1 juss
     90 just
      3 justera
      2 justerad
      4 justeras
      1 justerbar
      1 justerbara
      2 justering
      1 justeringar
      1 justeringarna
      1 justeringen
      1 justeringstemperatur
      2 justin
      1 justine
      1 justus
      4 juvéderm
      1 juveler
      1 juvelerare
      2 juvenil
      4 juver
      1 juvertumör
      5 juvret
      1 juvrets
      1 juxtaglomerulära
      1 jv
      1 jyllands
     17 k
      1 [k]
      1 k�
      2 ka
      1 kabatzinn
      2 kabel
      1 kabelisoleringen
      4 kabeln
      3 kabelprovare
      1 kabergolin
      1 kabi
      4 kablar
      1 kabylernas
      1 kackerlacka
      3 kad
      4 kadaver
      2 kadavret
      1 kadavrets
      1 kadinga
      1 kadmeia
     22 kadmium
      1 kadmiumabsorptionen
      1 kadmiumet
      1 kadmiummineral
      1 kadmiumupptaget
      1 kadmiumutsläppen
      1 kaducén
      1 kaféer
      4 kaffa
     15 kaffe
      1 kaffefärgad
      1 kaffein
      1 kaffekanna
      4 kaffelavemang
      1 kaffeplantager
      1 kaffeplantans
      1 kaffet
      1 kägelsnäckor
      3 kahunpapyrusen
      2 kairo
      2 kaj
      1 kajakpaddling
      1 kajal
      1 kajaleyeliner
      1 kajsamia
      2 käk
      1 kakao
      1 kakaobönan
      1 kakaobönor
      1 kakaohalt
      1 kakaohalten
      1 kakaolik
      3 käkar
      5 käkarna
      1 käkben
      1 käkbenet
      3 käke
      3 kakel
      1 kakelfix
      1 kakelfogar
      4 käken
      3 käkens
      3 kakexi
      1 käkinfektioner
      1 käkkirurg
      1 käkkirurger
      1 käkkirurgi
      1 käkkirurgiska
      1 kakko
      1 käkled
      1 käkleden
      1 käkleder
      1 käklederna
      1 käkmuskler
      1 käkmuskulatur
      2 käkmuskulaturen
      1 käkområdet
      1 kakor
      1 kakos
      1 kakosmi
      1 käkparti
      1 käksystem
     11 kal
      4 kål
      4 kala
      1 kalals
      1 kalanchoe
      1 kålblad
      1 kålbladen
      1 kålbladskompresser
      1 kalcifierade
      1 kalcifieras
      1 kalcifierat
      1 kalcineras
      2 kalcinering
      9 kalcitonin
      1 kalcitoninnivåer
     24 kalcium
      1 kalciumapatit
      1 kalciumbrist
      1 kalciumcitrat
      1 kalciumföreningar
      1 kalciumföreningarna
      1 kalciumfosfat
      2 kalciumhalt
      1 kalciumhalten
      1 kalciumhomeostas
      6 kalciumhydroxid
      7 kalciumhypoklorit
      1 kalciuminnehåll
      7 kalciumjoner
      1 kalciumjonerna
      1 kalciumkanaler
      1 kalciumkanalerna
     15 kalciumkarbonat
      1 kalciumkarbonatapatit
      1 kalciumkarbonatet
      5 kalciumklorid
      2 kalciumkloridhypoklorit
      1 kalciumnivå
      1 kalciumnivåerna
      1 kalciumomsättningen
      1 kalciumoxalat
      8 kalciumoxid
      1 kalciumpyrofosfatdihydrat
      2 kalciumsalter
      1 kalciumstearat
      1 kalciumsten
      2 kalciumstenar
      1 kalciumsulfat
      1 kalciumupptag
      1 kalciumutsöndring
      1 kalckar
      2 kalebasser
      1 kalebassvattenpipor
      2 kalender
      1 kålhuvudet
      1 kali
      1 kaliber
      1 kalibrerade
      1 kalifat
      1 kalifen
     11 kalifornien
      1 kaliforniens
      1 kalii
      1 kalilut
      1 kalinox
      2 kalippermetoden
     13 kalium
      1 kaliumaluminiumsulfat
      1 kaliumbikarbonat
      5 kaliumbromid
      3 kaliumcyanid
      1 kaliumcyaniden
      1 kaliumet
      1 kaliumgradient
      4 kaliumhydroxid
      1 kaliumhypoklorit
      1 kaliumjodat
     12 kaliumjodid
     12 kaliumjoner
      2 kaliumkarbonat
      1 kaliumklorid
      1 kaliumkloriden
      1 kaliumnitrat
      6 kaliumpermanganat
      2 kaliumsalter
      1 kaliumsåpa
      1 kaliumsåpor
      1 kaliumstegring
      1 kaliumsulfat
      1 kaliumvätesulfat
     12 kalk
      1 kalkaneussporre
      1 kalkartad
      1 kalkbildningen
      1 kalkblad
      1 kalkbladen
      2 kalken
      1 kalkfattig
      3 kalkhorn
      1 kalkkvävemetoden
      2 kalkrik
      1 kalkspat
      7 kalksten
      1 kalkyl
      9 kall
     20 kalla
     18 källa
      1 [källa
    292 kallad
    245 kallade
     70 kallades
      1 källafiltermodellen
     15 källan
      1 kallande
      1 källans
     22 kallar
      5 kallare
      2 källare
    813 kallas
      1 kallasläktet
    128 kallat
     11 kallats
      2 kallaväxter
      2 kallblodiga
      1 kallblodigt
      5 kallbrand
      1 kallde
      1 kalle
      2 kallelse
      1 källenius�svenson
      1 källkod
      1 kallmangel
      1 kallmanglar
      2 kallmanns
      2 källmaterialet
      1 kallmurade
      1 kallnat
      1 kallocain
      1 kallor
     64 källor
      1 källorna
      1 kallpressning
      1 kallrökta
      1 kallsläktet
      1 källsorteras
      1 kallsvetsning
      2 kallsvett
      1 kallsvettig
      1 kallsvettning
      1 kallsvettningar
     22 kallt
      1 kallvatten
      1 kallvattenkuranstalter
      1 kallvattenkuren
      5 kalmar
      1 kalmartrakten
      3 kalorier
      3 kaloriintag
      1 kalotypitekniken
      1 kålrötter
      1 kålsläktet
      1 kalsoho
      1 kalsonger
      1 kålsortertill
      3 kalv
      3 kalvar
      1 kalvarna
      1 kalvmage
      1 kalvmärkningstiden
      3 kam
      1 kamel
      2 kameldjur
      2 kamen
      8 kamera
      2 kameran
      1 kameror
      6 kamfer
      1 kamferartad
      2 kamfersyra
      1 kami
      1 kamikazeattackerna
      1 kaminireaktorerna
      1 kamliknande
      1 kammar
     29 kammare
      6 kammaren
      2 kammarens
      3 kammarflimmer
      1 kammarklaffarna
      1 kammarmusik
      3 kammarrätten
      1 kammarrättens
      1 kammarstängningarna
      1 kammarvätskan
      1 kammarvattnet
      1 kammens
      1 kammer
      1 kammre
      1 kamning
      1 kamomillextrakt
      2 kamouflage
      1 kamouflagefärger
      1 kamov
      4 kamp
      3 kämpa
      1 kämpade
      3 kampanj
      4 kampanjen
      3 kampanjer
      1 kämpar
      1 kämpat
      1 kämpe
      4 kampen
      1 kampmötena
      3 kampo
      1 kamporecept
      2 kamprespons
      1 kampresponsen
      2 kampsporter
      2 kampsportsskolor
      1 kamrar
     11 kamrarna
      2 kamrarnas
      3 kamrat
      4 kamrater
      1 kamratföreningar
      1 kamratrelationer
      1 kamratstöd
      1 kamskivling
   7701 kan
     34 kanada
      1 kanadafläder
      1 kanadas
      4 kanadensiska
      1 kanadensiske
      1 kanadensiskfödde
     10 kanal
      4 kanalen
     12 kanaler
      1 kanalerna
      1 kanalisera
      1 kancer
    100 känd
    144 kända
      1 kandahar
     11 kände
      2 kandidat
      1 kandidaten
      1 kandidater
      6 kandidatexamen
      1 kandidatgener
      2 kandidatprogrammet
      1 kandidera
      1 kandidos
      1 kändis
      3 kändisar
      1 kändisars
      1 kändisen
      1 kandy
      1 kanebo
      2 kanel
      1 kängor
      3 kängurumetoden
      1 kanin
      6 kaniner
      2 kanji
      1 kankunde
     91 känna
      1 kannan
      2 kännande
     21 kännas
      1 kännbar
      3 kännbara
      1 kannbrosk
      2 kannbrosken
      1 kannbroskens
      1 kannbroskkannbroskmuskeln
      7 kännedom
      1 kanner
    132 känner
      2 kanners
      1 kännetäcken
      1 känneteckande
     32 kännetecken
      1 kännetecknad
      7 kännetecknande
      1 kännetecknandes
     14 kännetecknar
     57 kännetecknas
      3 kännetecknet
      2 kannibalism
      1 kannibalistiska
     31 känns
      1 kanoniska
      2 kansas
      1 kansasii
     12 känsel
      5 känselbortfall
      2 känselcell
      2 känselförlust
      1 känselförlusten
      1 känselintryck
      5 känseln
      1 känselnedsättning
      1 känselnerverna
      1 känselplattor
      1 känselrubbningar
      3 känselspröt
      1 känselstörningar
     69 kanske
     69 känsla
     28 känslan
     27 känslig
     39 känsliga
      9 känsligare
      4 känsligast
      1 känsligaste
     33 känslighet
     14 känsligheten
      1 känsligheter
      1 känsligsom
      8 känsligt
      1 kanslist
      2 känslo
      1 känslobortfall
      1 känsloladdade
      2 känsloliv
      4 känslolivet
     17 känslomässig
     18 känslomässiga
     12 känslomässigt
     89 känslor
      1 känsloreaktioner
      1 känsloreglerande
      4 känslorna
      1 känslorörelse
      1 känslosamhet
      1 känslosamme
      1 känslostrukturerna
      1 känslosvängningar
      3 känslotillstånd
      1 känsloupplevelser
      1 känsloutbrott
      1 känslovärld
     21 kant
     89 känt
      1 kantad
      1 kantagonist
      1 kantar
      1 kantas
      9 kanten
      7 kanter
      5 kanterna
      1 kantiga
      1 kantigt
      1 kantnerver
      1 kantnerverna
      1 kanton
      1 kants
      3 känts
      1 kantvinklar
     12 kanyl
      6 kanylen
      1 kanylens
     11 kanyler
      1 kanylerad
      1 kanyls
      6 kaos
      1 kaotiska
      2 kaotiskt
      9 kap
      1 kåpa
      6 kapabel
      1 kapabla
      1 kapacitans
      2 kapacitansen
     16 kapacitet
      3 kapaciteten
      1 kapad
      1 kåpan
      2 kapas
      1 kapats
      2 kapell
      1 kapellvred
      1 kapha
      2 kapillär
      1 kapillära
      1 kapillärbädd
      1 kapillärbädden
      1 kapillärblod
      9 kapillären
      1 kapillärens
     21 kapillärer
     13 kapillärerna
      1 kapillärernas
      1 kapillärnätet
      2 kapillärsystem
      1 kapillärsystemet
      1 kapillärt
      1 kapillärtryck
      2 kapillärtrycket
      1 kapillärväggar
      1 kapillärväggen
      1 kapitalisten
      1 kapitalt
      8 kapitel
      1 kaplan
      1 kapnograf
      4 kaposis
      2 käpp
      2 kappadokien
      4 käppar
      1 käpparna
      3 käppen
      1 kapprustning
      1 käpptekniken
      1 kapris
      1 kaprolakton
     10 kapsel
      2 kapselendoskopi
      1 kapselendoskopin
      1 kapseltänder
      1 kapsla
      1 kapslad
      6 kapslar
      1 kapslas
      1 kapsling
      1 kapsomerer
      1 kapstaden
      3 kapsulotomi
      1 kapsutolomi
      1 kapten
      1 kaptenen
      5 kär
      2 kära
     31 karaktär
      5 karaktären
      7 karaktärer
      1 karaktärernas
      1 karaktäriserad
      1 karaktäriserar
     11 karaktäriseras
      1 karaktäriserat
      1 karaktariskt
      2 karaktäristika
      4 karaktäristisk
      4 karaktäristiska
      6 karaktäristiskt
      5 karaktärsdrag
      2 karaktärsdragen
      1 karaktärsfel
      1 karaktärsfullt
      1 karaktärsneuros
      1 karaktärsneuroser
      3 karakterisera
      1 karakteriserade
      1 karakteriserar
     16 karakteriseras
      2 karakteriserat
      1 karakterisering
      2 karakteristika
     11 karakteristisk
     10 karakteristiska
      4 karakteristiskt
      1 karäkteristiskt
      1 karamoja
      1 karankawaindianerna
     13 karantän
      1 karantänsanstalt
      1 karantänsperioder
      2 karat
      1 karavaner
      1 karbad
      1 karbamat
      2 karbamazepin
      1 karbamazepinbaserade
      2 karbamidperoxid
      4 karbaminohemoglobin
      1 karbaminohemoglobinet
      6 karbapenemer
      1 karbin
      1 karbolchampinjon
      2 karbolsyra
      1 karbonat
      1 karbonatapatit
      1 karbonylgrupp
      1 karboxihemoglobin
      3 karboxylgrupp
      1 karboxylgrupperna
      5 karboxylsyra
      3 karboxylsyror
      2 karbunklar
      2 karcinoid
      1 karcinoida
      1 karcinoider
      1 karcinoidsyndrom
      1 karcinom
      1 kardia
      1 kardinalsaft
      1 kardinalsafternas
      4 kardinalsymtom
      1 kardinalsymtomet
      2 kardioacceleratoriska
      1 kardiogen
      1 kardiolog
      5 kardiologer
      4 kardiologi
      2 kardiomyopati
      1 kardiomyopatier
      5 kardiovaskulär
      7 kardiovaskulära
      1 kardiovaskul�r
      1 kareler
      1 karelsk
      1 karelska
      1 karensregler
      1 kårer
      1 karettsköldpadda
      1 karettsköldpaddorna
      6 kärfve
      2 karibien
      8 karies
      1 kariesaktivitet
      2 kariesangrepp
      2 kariesangreppen
      1 kariesorsakande
      1 kariesprovocerande
      1 kariesuppkommande
      4 karin
      1 käringknut
      1 karisma
      1 karjakin
     17 karl
     33 kärl
      1 kärlavledning
      1 kärlavslappande
      1 karlaxel
      1 kärlbiten
     19 kärlek
      3 kärleken
      1 kärleksäpplen
      1 kärleksbehov
      1 kärleksberoende
      1 kärleksfattiga
      1 kärleksfull
      1 kärlekshormon
      1 kärleksrelation
      4 kärleksrelationer
     14 kärlen
      1 karlén
      1 kärlens
      1 karlerik
     14 kärlet
      2 kärlets
      1 kärlförlängning
      1 kärlformade
      1 kärlförträngningarna
      1 kärlförträngningarnas
      1 karlgustav
      1 kärlinflammation
      1 kärlkirurgi
      9 kärlkramp
      1 kärllumen
      1 kärlmissbildning
      1 kärlmissbildningar
      1 kärlnät
      1 kärlresistans
      1 kärlresistansen
      1 kärlrespons
      5 kärlsammandragande
      1 karlsbadersalt
      1 karlsbadervatten
      1 kärlsektionen
      5 kärlsjukdom
     14 kärlsjukdomar
      1 kärlsjukdomen
      1 kärlskada
      1 karlskrona
      3 kärlsonografi
      1 karlstad
      1 kärlstrukturer
      1 kärlsystem
      1 kärlsystemet
      1 kärltillväxten
      1 kärlträdet
      1 kärlvägg
      7 kärlväggarna
     12 kärlväggen
      1 kärlväxt
      1 kärlvidgning
      1 karma
      1 karmalagen
      1 karmar
      1 karmayoga
      1 kärmehinen
      1 kärmet
      9 kärna
      7 kärnan
      2 kärnans
      3 kärnbränsle
      1 kärndna
      1 karnevalen
      1 kärnfasväxling
      1 kärnfrågan
      1 kärnklyvning
      2 kärnkraft
      1 kärnkraftsindustri
      1 kärnkraftsolycka
      1 kärnkraftsprogram
      3 kärnkraftverk
      1 kärnladdningar
      1 kärnmaterial
      7 kärnor
      1 kärnorna
      1 kärnreaktor
      5 kärnreaktorer
      1 kärnreceptorer
      1 kärnsprängningarna
      1 kärnupplevelse
      9 kärnvapen
      2 kärnvapenprogrammet
      1 karofyter
      1 karolina
     38 karolinska
      1 karotenoiden
      1 karotenoider
      1 karotisblodkärlet
      1 karotyper
      2 karpaltunneln
      1 karpaltunnelns
      9 karpaltunnelsyndrom
      1 karpaltunnelsyndromär
      1 karpeller
      1 karpos
      1 karposis
      1 kärr
      7 karragenan
      1 karragentång
      4 karriär
      1 karsianus
      1 kartageners
      1 kartfjäril
      1 karthagiske
      1 kartlade
      3 kartlades
      8 kartlägga
      5 kartlägger
      5 kartläggning
      1 kartläggningen
      2 kartlagt
      1 kartlagts
      1 kartong
      1 kartor
      1 karusell
      1 karvakrol
      1 karvinskianus
      1 karyotyp
      3 kasam
      1 kaseös
      1 kasinot
      1 kasjunöt
      2 kaskad
      1 kaspiska
      2 kassava
      3 kasseras
      1 kasserats
      1 kassettband
      1 kassettfilter
      1 kassor
      1 kassunarbetarna
      2 kassunen
      1 kassuner
      3 kast
     10 kasta
      1 kastade
      1 kastanjenötter
      7 kastar
      6 kastas
      1 kastmaskiner
      1 kastning
      3 kastration
      1 kastratsångare
      1 kastrera
      2 kastrerade
      1 kastrerades
      2 kastrerat
      6 kastrering
      2 kastrull
      1 kastruller
      1 kastväsendet
      1 kat
      2 katabol
      1 katabola
      1 kataktärsneurotiska
      4 katalas
      1 katalasnegativa
      7 katalepsi
      1 katalepsiattack
      2 katalog
      1 kataloger
     13 katalysator
      1 katalysera
      8 katalyserar
      3 katalyseras
      1 katalyserat
      3 katalytisk
      1 katalytiska
      1 katalytiskt
      1 katameniell
      1 katameniella
     10 kataplexi
      2 kataplexiattackerna
      5 kataplexin
      1 kataplexis
      1 katapultstol
      4 katarakt
      1 kataraktkirurgi
      1 katarina
      1 katarr
      7 katastrof
      1 katastrofala
      1 katastrofalt
      2 katastrofartad
      3 katastrofen
      9 katastrofer
      3 katastrofmedicin
      1 katastrofplats
      1 katastrofplatser
      2 katastroftankar
      1 katastroftanken
     12 kataton
      1 katatona
     11 katatoni
      2 katatont
     10 katatreni
      1 katatrenin
      1 katatrenipatienter
      2 kate
     18 kategori
     26 kategorier
      3 kategorierna
     11 kategorin
      3 kategorisera
      2 kategoriserade
      2 kategoriserar
     10 kategoriseras
      2 kategorisering
      1 kategoriseringen
      1 kategorisk
      2 katekol
      8 katekolaminer
      1 katekolaminerna
      1 katekolometyltransferas
      1 kateogorin
     24 kateter
      1 kateterar
      1 kateterbehandling
      1 kateterformat
      7 kateterisering
      1 kateteriseringen
      1 kateterlängden
     13 katetern
      1 kateterspetsen
      1 kateterteknik
      1 kateterundersökning
     15 katetrar
      2 katetrarna
      2 katetrisering
      1 katharsis
      1 kåthet
      1 kathon
      1 katie
      1 katin
      3 katinon
      1 katinonfamiljen
      1 katjon
      1 katjonaktiva
      1 katjoner
      1 katod
      1 katoden
      1 katodstråleoscillograf
      1 katodstråleoscilloskopen
      1 katodstrålerör
      5 katodstråleröret
      2 katoliker
      9 katolska
      1 katrineholm
     11 katt
      1 kattan
      3 kattavföring
      3 kattdjur
      7 katten
      3 kattens
     32 katter
      3 kätteri
      2 katterna
      1 katters
      1 kattgut
      1 katthår
      4 kattlådan
      1 kattöga
      1 kattögereflexen
      1 kattorganisationer
      1 kattorganisationerna
      1 kattparasit
      1 kattraser
      1 katttarm
      1 kattuggla
      2 kattungar
      1 kaudalt
      1 kaukasier
      1 kaukasisk
      8 kaukasus
      2 kaulitz
      2 kausal
      1 kausala
      2 kausalitet
      3 kausalt
      1 kauteri
      1 kauterisering
      2 kavelbräden
      2 kaviteten
      2 kaviteterna
      1 kaxinawa
      1 kayanfolket
      1 kazakhstan
      1 kazakstan
      1 kazdin
      1 kazonogla
      1 kbk
     25 kbt
      1 kbtbaserad
      1 kbtterapi
      5 kcal
      1 kcn
      1 kcnj
      2 kda
      1 keats
      6 kedja
      9 kedjan
      2 kedjereaktion
      1 kedjereaktionen
      1 kedjeröker
      2 kedjetransplantation
      7 kedjor
      1 kees
      1 kefale
      1 kegel
      1 kegelträning
      1 keiron
      2 keith
      1 keiths
      1 kejsar
      1 kejsare
      3 kejsaren
      1 kejsarens
      1 kejsarinnan
     42 kejsarsnitt
      1 kejsarsnittens
      5 kejsarsnittet
      1 kejsarsnittsandel
      1 kejsarsnittsfrekvens
      1 kejsarsnittsfrekvensen
      1 kelade
      1 kelidon
      2 keller
      1 kells
      1 keloid
      1 kelsos
      1 keltisk
     22 kemi
      1 kemiföretaget
      4 kemikalie
      1 kemikalieexport
      1 kemikalieexportförbud
      1 kemikaliefrisättning
      3 kemikalieindustrin
      1 kemikalieindustris
      5 kemikalieinspektionen
      1 kemikalielagstiftning
      1 kemikaliemyndighet
      3 kemikaliemyndigheten
      3 kemikalien
      1 kemikalieproducenter
      1 kemikalieproducenterna
      1 kemikalieproduktionen
     47 kemikalier
      4 kemikalierna
      2 kemikaliers
      1 kemikalietillverkarna
      5 kemin
      1 kemins
      1 kemira
      1 kemishowexperiment
     67 kemisk
     96 kemiska
     26 kemiskt
      1 kemispråk
     16 kemisten
      3 kemister
      1 kemisterna
      1 kemodestruktiv
      1 kemokiner
      2 kemomekanisk
      1 kemoreceptor
      7 kemoreceptorer
      8 kemoreceptorerna
      1 kemoreduktion
      1 kemoterapeutisk
      1 kemoterapeutiskt
     14 kemoterapi
      1 kemtvättas
      1 kemtvättautomater
      3 kennedy
      1 kennel
      5 kennelhosta
      1 kennelklubben
      1 kennlar
      1 kenofobi
      3 kent
      1 kentauren
      2 kentucky
      3 kenya
      1 kephal�
      1 kephal�huvud
      1 kepoxidreduktas
      1 keramik
      1 keramiska
      2 keramiskt
      1 keratinas
      2 keratinet
      1 keratinfibriller
      3 keratit
      1 keratitis
      1 kermeinen
      3 kermesbär
      4 kernigs
      1 kerry
      1 kerstin
      4 kes
      3 ketamin
      1 ketchupeffekt
      1 keto
      7 ketoacidos
      1 ketobemidon
      1 ketogan
      2 ketogen
      1 ketoglukonsyra
      1 ketogruppen
      1 ketokropparnas
      5 keton
      7 ketoner
      1 ketonerna
      7 ketonkroppar
      1 ketonkropparna
      1 ketonkroppsbildning
      1 ketonproduktionen
      5 ketonsyraförgiftning
      1 ketonvärden
      8 ketos
      1 ketosbildningen
      1 ketosis
      1 ketosyra
      4 kev
      1 kevlarmaterial
      1 kex
      2 key
      1 kfiskada
      1 kfs
      1 kfs]
     37 kg
      1 �kg
      1 kgb
      4 kgm
      1 kg�min
      2 kh
      1 kha
      1 khan
      1 khnum
      3 khz
      7 ki
      1 kiai
      1 kiba
      6 kick
      3 kicken
      1 kidnapparenkidnapparna
      2 kidnapparna
      1 kidnappning
      1 kidnappningsoffer
      1 kiedis
      2 kiel
      1 kiels
      1 kiflöde
      1 kifs
      1 kikärter
     21 kikhosta
      1 kikhostebakterier
      1 kikhosteliknande
      1 kikhostesmitta
      1 kikhostliknande
      1 kikhoststadiet
      1 kikningarna
      2 kilar
      1 kilbenet
      1 kille
      1 killed
      1 killian
      2 killing
     23 kilo
     11 kilogram
      1 kilokalorier
      2 kilometer
      2 kilometers
      1 kilon
      1 kilovolt
      1 kilskrifter
      1 kimssi
     60 kina
      2 kinas
      2 kinasdomänen
      2 kinase
      1 kinashämmare
      1 kinasyra
      2 kind
      3 kinder
      3 kinderna
      1 kindesalter
      1 kindtänderna
      1 kinematiska
      3 kineret
      2 kineser
      1 kineserna
      2 kinesernas
      1 kinesiologer
      3 kinesiologi
      1 kinesiologin
      1 kinesis
     12 kinesisk
     16 kinesiska
      1 kinetik
      1 kinetiska
      3 king
      6 kinin
      1 kininallergi
      1 kininet
      2 kinolonen
      8 kinoloner
      1 kinolonerna
      1 kinolonresistens
      1 kinsey
      1 kiptjakkhanen
      2 kiral
      1 kirlianfotografering
     17 kiropraktik
     10 kiropraktiken
      3 kiropraktikens
      1 kiropraktikskolor
      7 kiropraktisk
      3 kiropraktiska
      8 kiropraktor
      1 kiropraktorbildningen
     14 kiropraktorer
      1 kiropraktorerna
      1 kiropraktorernas
      3 kiropraktorers
      3 kiropraktorhögskolan
      1 kiropraktorn
      1 kiropraktorutbildning
      1 kiropraktorutbildningar
      2 kiropraktorutbildningen
      1 kirskål
      6 kirurg
      1 kirurgavdelningen
     14 kirurgen
     11 kirurger
      4 kirurgerna
      1 kirurgernas
    109 kirurgi
      1 kirurgie
      1 kirurgimetoder
      7 kirurgin
      4 kirurgins
     52 kirurgisk
     50 kirurgiska
     52 kirurgiskt
      1 kirurgknut
      1 kirurgläkare
      1 kiseldioxid
      1 kiseldioxidyta
      1 kiselgur
      2 kiselpulver
      1 kiselpulvret
      1 kiselsanering
      1 kiseru
      1 kiseruer
      2 kiserun
      1 kiske
      9 kissa
      1 kissande
      3 kissar
      1 kisseflaska
      1 kissing
      1 kisslarm
      1 kisspeptin
      2 kista
      1 kitazato
      1 kitsune
      1 kittfärgad
      2 kittlande
      1 kittlar
      1 kittlas
      1 kiurgiskt
      1 kiva
      1 kiwiavokado
      1 kiyoshi
      1 kj
      2 kjell
      1 kjolarna
      1 kjolen
      1 kjonkanaler
      5 kl
      1 klä
      1 kläckas
      1 kläckning
      2 kläckningen
      1 kläckningsplatser
     14 kläcks
      4 kläcktes
     48 klåda
      8 klådan
      1 klådavanligen
      1 kladd
      1 klädd
      1 kladda
      7 klädda
      1 klåddämpande
      1 kladdar
      2 klädde
      2 kläddes
      2 kladdiga
      1 klädedräkt
      1 klädedräkten
     54 kläder
     10 kläderna
      1 klädernapälsen
      6 klädesplagg
      1 klädfrihet
      1 klådfritt
      2 klädhängare
      1 klädhängaren
      1 klädklämma
      2 klädkod
      1 klädkoder
      1 klådlindrande
      1 klädlinjen
      1 klädlöss
      1 klädnad
      2 klädnypa
      2 klädnypan
      3 klädnypor
      1 klädnyporna
      2 kladogram
      1 klädproduktionen
      4 klädsel
      1 klädseln
      4 klädstreck
      3 klädstrecket
      1 klädtvätt
      1 klädvaruhuset
      1 klaffande
      5 klaffar
      7 klaffarna
      1 klaffarnas
      1 klaffsjukdomar
      1 klaga
      1 klagade
      1 klagande
      1 klagar
      2 klagomål
      1 klagomålen
      4 kläm
      1 klämflaska
      8 klämma
      1 klämmare
      1 klammer
      3 klämmer
      3 kläms
     13 klamydia
      1 klamydiadiagnoser
      2 klamydiainfektion
      1 klamydiaprov
      1 klamydiase
      1 klamydiasmitta
      1 klamydiasmittade
      3 klamydiatest
      1 klamydiatestnu
      1 klamydiavarianten
      3 klander
      1 klandrar
      1 klandrats
      3 klang
      2 klänga
      1 klängande
      3 klänge
      1 klängen
      1 klängena
      1 klänger
      1 klangfärgen
      1 klänning
      1 klänningar
      1 klänningsliknande
      2 klappa
      1 klappade
      2 klappar
      1 klapphingstar
      1 klaproth
     23 klar
      1 klär
     43 klara
      3 klarade
     51 klarar
      4 klarat
      1 klarcellscarcinom
      1 klardröm
      1 klardrömmande
      3 klardrömmar
      3 klargjorde
      1 klargör
      4 klargöra
      1 klargörande
      1 klargörs
      1 klarlades
      7 klarlagd
      2 klarlagda
      2 klarlägga
     15 klarlagt
      1 klarnat
      1 klarningsmedel
      1 klarröd
      1 klarröda
      1 klarrött
     24 klart
      1 klartext
      1 kläs
      6 klasar
      4 klase
     17 klass
      1 klassad
      2 klassade
      3 klassades
      1 klassar
     31 klassas
      4 klassat
      1 klassats
     12 klassen
     12 klasser
      4 klasserna
     10 klassificera
      1 klassificerade
      1 klassificerades
      2 klassificerar
     29 klassificeras
      1 klassificerat
      2 klassificerats
     20 klassificering
      8 klassificeringen
      2 klassificeringssystem
      1 klassificieras
     14 klassifikation
      1 klassifikationen
      1 klassifikationerna
      1 klassifikationssystem
      1 klassifikationssystemet
      3 klassifikationstest
      2 klassiker
      1 klassindelning
     36 klassisk
     36 klassiska
      4 klassiskt
      1 klassning
      1 klasstillhörighet
      1 klatschandet
      1 klatskins
      3 klätt
      3 klätten
      4 klättersumak
      4 klättra
      3 klättrande
      3 klättrar
      1 klättrare
      1 klättrat
      1 klättring
      1 klätts
      1 klaus
      4 klaustrofobi
      1 klebs
      7 klebsiella
      4 klein
      1 klen
      4 kleopatra
      1 klepto
      1 kleptofili
      1 kleptoman
      1 kleptomaner
      9 kleptomani
      7 klia
      5 kliande
      1 kliandet
     11 kliar
      2 klibba
      2 klibbar
      1 klibbig
      2 klibbiga
      1 klibbighet
      3 klibbigt
      1 klibbnattskatta
      1 klichémässigt
      3 klick
      1 klickljud
      1 klient
      1 klientcentrerade
      1 klientcentrerat
     17 klienten
      7 klientenpatienten
      4 klientens
      5 klienter
      1 klienterna
      1 klienternas
      1 klienterpatienter
      3 klimakteriebesvär
      1 klimakteriebevärd
     23 klimakteriet
      4 klimakterium
     20 klimat
      5 klimatet
      1 klimatförändringar
      1 klimatförändringarna
      1 klimatförändringarnas
      1 klimatförändringen
      1 klimatförhållanden
      1 klimatkatastrofer
      1 klimatologiska
      1 klimax
      4 klindamycin
      1 kline
      2 klinefelters
      1 kling
      1 klinga
      1 klingande
      4 klingar
      2 klingbergs
      1 klingenberg
      8 klinik
      1 klinikblekning
      1 klinikchefsarbete
     16 kliniken
     11 kliniker
      8 klinikerna
      1 kliniks
     68 klinisk
     86 kliniska
      1 klinisk�medicinska
     34 kliniskt
      1 klinken
      1 klinker
      1 klinkik
      3 klippa
      2 klippas
      1 klippavsats
      1 klippdel
      1 klippel
      1 klippelfeils
      5 klippeltrenaunay
      1 klippeltrénaunay
      2 klippeltrenaunays
      2 klippiga
      2 klippning
      1 klippta
      1 klipptes
      1 klippts
      1 klisterfläckar
      2 klisterremsa
      1 klistrad
      1 klistrar
      4 klistras
     15 klitoris
      1 klitorism
      1 klitorispiercing
      1 klitoristoppen
      2 klitoromegali
      1 klivit
      1 klo
      1 kloakdjur
      1 kloaker
      2 kloaköppning
      9 klocka
      3 klockan
      5 klockformade
      1 klockjulros
      1 klocklik
      2 klocklika
      1 klockliljesläktet
      2 klockor
      1 klockorna
      1 klockrike
      1 klockringningar
      1 klockslag
      1 klockslager
      1 klocktest
      3 klok
      4 kloka
      1 klokt
      1 kloliknande
      1 klomipramin
      4 klon
      1 klonal
      3 klonen
      1 kloner
      1 klonselektionsteorin
      3 klonus
      1 klopidogrel
     28 klor
      2 klorakne
      2 kloralhydrat
      2 kloramfenikol
      1 kloranil
      1 kloratomer
      1 klorattillverkning
      2 klorbaserade
      1 klorbensen
      1 klorbensenetan
      1 klorblekning
      1 klordesinfektion
      1 klordesinfiktion
      1 klordiklorfenoxifenol
      7 klordioxid
      1 klordioxiden
      3 klorerade
      2 kloreras
      2 klorering
      7 kloretan
      1 kloretanol
      1 klorex
      1 klorfenol
     11 klorgas
      6 klorhexidin
      1 klorhexidinpreparat
      3 klorid
      1 kloriden
      1 kloridjoner
      1 kloridkanaler
      4 klorin
      1 klorjoner
      7 klorkalk
      1 klorlukt
      1 klorluktande
     11 klormetan
      1 klormetanföreningar
      1 klormezanon
      1 klorna
      1 kloroamfenikol
     26 kloroform
      2 kloroformanestesi
      2 kloroformliknande
      1 kloroforms
      2 klorofyll
      1 klorokin
      3 kloster
      1 klosterträdgårdarna
      2 klostren
      1 klot
      1 klotrund
      1 klotrunda
      1 klotsar
      1 klovård
      2 klövarna
      1 klövbärande
      1 klövhornet
      1 klövklipp
      1 klövsjuka
      1 klövspalten
      1 klövspaltseksem
      1 kloxacillin
      1 klozapin
      4 klubb
      3 klubbar
      1 klubbarna
      2 klubben
      1 klubbhus
      1 klubblag
      2 klubbyte
      3 klump
      2 klumpa
     10 klumpar
      1 klumparna
      1 klumpförebyggande
      3 klumpfot
      1 klumpfotliknande
      1 klumpkänsla
      1 klumprot
      1 klumprotsjuka
      3 klungor
      1 klusil
     10 klusiler
      1 klusiltypen
      1 klusiltyper
      9 kluster
      1 klustret
      1 kluven
      1 kluvet
      4 klyka
      1 klypa
      1 klysma
      1 klyva
      1 klyvbart
      2 klyver
      1 klyvning
      1 klyvningsprodukt
      4 klyvs
      5 km
      8 kmh
      1 �kmh
      1 kmno
      2 kmt
      2 kmtim
      1 kmtimme
     10 knä
      1 knacka
      1 knackar
      1 knackningar
      2 knåda
      1 knådas
      3 knådning
      1 knådningar
      2 knäet
      2 knäleden
      1 knäledens
      2 knäleder
      1 knälederna
      2 knäledsartros
      1 knäledsdysplasi
      7 knän
      7 knäna
      5 knapp
      3 knappar
      1 knappas
     13 knappast
      2 knappen
      1 knäpper
      2 knapphändig
      2 knäppningar
     28 knappt
      1 knapptryckande
      1 knapptryckning
      1 knarkfabriker
      2 knarr
      2 knarrande
      2 knarren
      1 knarrig
      1 knäskada
      1 knäskador
      1 knäskålen
      2 knäsvaghet
      7 knät
      1 knäts
      1 knick
      1 knipövning
      1 knipövningar
      1 knippe
      3 knippen
      4 kniv
      3 knivar
      1 knivblad
      1 knivens
      1 knivkastning
      2 knivlagen
      1 knivliknande
      1 knivslida
      1 knivsta
      1 knogarna
     14 knöl
     10 knölar
      3 knölarna
      3 knölen
      1 knölformad
      1 knölformig
      1 knöligt
      1 knölpåkar
      1 knopp
      1 knoppar
      2 knoppas
      2 knoppen
      1 knossospalatset
      1 knöt
      1 knotor
      2 knott
      1 knotten
      1 knottrig
      2 knottriga
      1 knottrighet
      9 knottror
      1 knowledge
      1 knox
      1 kns
      1 knubbiga
      1 knubbsälar
      1 knud
      1 knuff
      1 knuffa
      1 knuffade
      7 knut
      1 knuta
      2 knutar
     13 knuten
      8 knutet
      5 knutna
      4 knutor
      1 knutpunkter
      7 knyta
      2 knytas
      8 knyter
      2 knytits
      3 knyts
      8 ko
      1 kö
      5 koagel
      1 koaglet
      1 koagulas
      1 koagulasnegativa
      7 koagulation
      3 koagulationen
      1 koagulationfaktorerna
      1 koagulationfaktorn
      2 koagulationsfaktor
      5 koagulationsfaktorer
      2 koagulationsfaktorerna
      1 koagulationsförloppen
      2 koagulationsförmåga
      3 koagulationsförmågan
      1 koagulationshämmande
      1 koagulationsinducerad
      2 koagulationsproteiner
      4 koagulationssystemet
      8 koagulera
      2 koagulerar
      3 koagulerat
      5 koagulering
      2 koaguleringen
      1 koaguleringsförmåga
      1 koaguleringsprocessen
      5 koalitionen
      1 koalitioner
      1 koanalatresi
      1 koanophyllon
      1 kobent
      1 kobenthet
      1 köbildning
      3 kobolt
      1 koboltkanonen
      1 kōbon
      1 kobra
      5 koch
      1 kock
      2 kockar
      1 kocken
      3 kocker
      1 kockhandduk
      2 kod
      1 koda
      1 kodaikanal
      2 kodak
      1 kodande
     11 kodar
      1 kodas
      3 kodein
      1 koder
      1 kodningen
      1 kodsystemet
      1 koeberlé
      1 koelia
      1 köer
      1 kofaktor
      1 kofaktorn
     30 koffein
      1 koffeinberoende
      1 koffeinet
      1 koffeinets
      1 koffeinförgiftning
      1 koffeinintag
      1 koffeinkällor
      1 koffeinkoncentration
      1 koffeinlösning
      4 kofferdam
      1 kofferdamduken
      1 kofferdamen
      1 kofi
      1 koger
      4 kognition
      4 kognitionen
      1 kognitions
      1 kognitionspsykologi
     69 kognitiv
     46 kognitiva
      7 kognitivt
      2 koh
      2 koherens
      1 kohorn
      2 kohort
      1 kohorter
      2 kohortstudie
      1 kohortstudier
      1 kohoul
      1 koiliakos
      4 kök
      6 koka
      1 kokad
      1 kokades
      9 kokain
      1 kokainets
      2 kokande
      1 kokapparat
      4 kokar
      2 kokard
      7 kokas
      1 köken
      5 köket
      1 kökets
      1 kokhett
      1 kokkärl
     12 kokning
      1 kokningen
      2 kokong
     13 kokoppor
      1 kokoppviruset
      1 kokos
      1 kokosmjölk
      1 kokosnötolja
      1 kokosnötter
      1 kokosolja
      5 kokpunkt
      1 koks
      7 koksalt
      5 koksaltlösning
      1 koksaltproteser
      1 kökshandduk
      1 kökshanddukar
      1 kökshandduken
      1 köksknivar
      1 köksluckor
      1 kökspapper
      2 köksredskap
      1 köksredskapen
      1 kökssläng
      1 köksspecialister
      1 koksverk
      1 kokt
      1 kokta
      1 kokvagnar
      1 kokvatten
     25 kol
      2 köl
      2 kola
      1 kolanalys
      1 kolangiocarcinom
      1 kolanöten
      1 kolarbetarlungor
     14 kolatom
      5 kolatomen
     14 kolatomer
      1 kolatomerna
      1 kolbe�schmitt
      8 kölbröst
      1 kolchicin
      2 koldifluorid
     68 koldioxid
      4 koldioxiden
      4 koldioxidens
      1 koldioxidfrisättning
      1 koldioxidgas
      1 koldioxidhalt
      3 koldioxidhalten
      1 koldioxidis
      1 koldioxidkoncentration
      1 koldioxidmolekyl
      1 koldioxidpartialtrycket
      1 koldioxidtrycket
      1 koldisulfid
      1 köldkänslighet
      1 köldmaskinerier
      3 köldmedium
      1 köldskada
      1 köldskadad
      4 köldskador
      1 köldtåliga
      1 kolecystokinin
      1 kolecystokininpankreozymin
      1 koledokus
      2 koleldade
     16 kolera
      2 kolerabakterien
      2 koleraepidemi
      1 koleraepidemier
      1 koleraepidemin
      1 kolerafall
      7 koleran
      1 kolerans
      1 kolestas
      1 kolestaslymfödemsyndrom
     19 kolesterol
      1 kolesterolabsorptionshämmaren
      2 kolesterolet
      1 kolesterolhalten
      1 kolesterolkoncentrationen
      1 kolesterolnivån
      1 kolesterolsänkande
      1 kolesterolvärdet
      1 kolet
      2 kolfiber
      1 kolfiberdetaljer
      1 kolfiltermattor
      2 kolföreningar
      1 kolförgasning
      4 kolhydrat
      1 kolhydratbrist
     40 kolhydrater
      1 kolhydraterenergi
      9 kolhydraterna
      1 kolhydraternas
      2 kolhydratfattig
      1 kolhydratfattiga
      1 kolhydratinnehåll
      5 kolhydratintag
      5 kolhydratintaget
      1 kolhydratkällan
      1 kolhydratkedjor
      1 kolhydratkonsumtion
      1 kolhydratrik
      3 kolhydratrika
      1 kolhydratsförsöket
      1 kolhydratsintaget
      1 kolhydratsorter
      1 kolibakterier
      1 koliforma
      4 kolik
      1 kolikliknande
      1 koliksmärtor
      1 kolin
      1 kolinerg
      4 kolinerga
      1 kolinesteras
      1 kolinesterashämmare
      1 kolingen
      2 kolingens
     15 kolit
      1 kolk
      5 kolkedja
      3 kolkedjan
      1 kolkedjedelen
      1 kolkedjor
      1 kolkicin
      3 koll
      3 kolla
     11 kollagen
      1 kollagenbaserad
      1 kollagenfiber
      1 kollagenfibrer
      1 kollagenfibrerna
      1 kollagenlager
      1 kollagenrik
      1 kollagenskikt
      1 kollagensyntesen
      4 kollaps
      1 kollapsa
      2 kollapsade
      1 kollapsat
      3 kollapsterapi
      1 kollar
      1 kollas
      1 kollateralkärl
      2 kollega
      1 kolleger
      8 kollegor
      1 kollekt
      1 kollektion
      2 kollektiva
      3 kollektivavtal
      2 kollektivistiska
      1 kollektivistiskt
      3 kollektivt
      1 kollektivtrafik
      2 kollektivtrafiken
      1 kollidera
      2 kolliderar
      2 kollimator
      1 kollimatorer
      1 kollimering
      3 kollision
      1 kollodiumprocesserna
      1 kollodiumtorrplåtar
      1 kollodiumvåtplåtar
      1 kolloidal
      1 kolloidosmatiska
      4 kolloidosmotiska
      1 kolloidosmotiskt
     26 kolmonoxid
      1 kolmonoxiden
      5 kolmonoxidförgiftning
      2 kölna
      8 kolobom
      2 kolobomet
      1 kolokvint
      4 kolon
      1 koloncancer
      4 koloni
      1 kolonial
      1 koloniala
      1 kolonialadministrationen
      1 kolonialisering
      1 kolonialväldet
      3 kolonibildande
      6 kolonier
      1 kolonisation
      1 kolonisationen
      1 kolonisationer
      1 kolonisatörer
      2 kolonisera
      4 koloniserade
      1 koloniserades
      4 koloniserar
      1 koloniserat
      1 koloniserats
      1 koloniseringen
      1 kolonistimulerande
      1 kolonivis
      1 kolonn
      2 kolonnen
      1 kolonnmetoder
      1 kolonnskaft
      2 kolorektal
      1 kolorektalkirugi
      1 kolos
      5 koloskopi
      3 kolostomi
      1 kolostomins
      3 kolostrum
      1 koloxid
      1 koloxidförgiftning
      1 kolstift
      4 kolstybb
      1 kolsva
      1 kolsvart
      1 kolsvavla
      1 kolsvavlelösning
      5 kolsyra
      1 kolsyrad
      1 kolsyran
      1 kolsyras
      1 kolsyrehaltigt
      1 kolt
      1 koltabletter
      2 koltåldern
      1 koltetraklorid
      1 kolumn
      1 kolumner
      2 kolv
      7 kolväte
      1 kolväteförening
      1 kolvätegrupp
      6 kolväten
      1 kolvätet
      1 kolväteutsläpp
      2 kölvatten
      2 kölvattnet
      1 kolven
    198 kom
     42 koma
      1 komaanfall
      1 komärket
      1 komarovii
      1 komatillståndet
      1 komatös
      1 komatöst
      1 kombattanter
      1 kombimodell
    136 kombination
     17 kombinationen
     13 kombinationer
      2 kombinationerna
      2 kombinationsbehandling
      2 kombinationspiller
      4 kombinationspreparat
      1 kombinationsschampon
      1 kombinationsvaccin
      1 kombinationsvaccinet
      9 kombinera
     12 kombinerad
      5 kombinerade
      4 kombinerades
      7 kombinerar
     34 kombineras
     13 kombinerat
      6 kombucha
      1 kombuchasvampen
      1 komdovaranen
      1 komedi
      8 komet
      1 kometmetoden
      6 komfort
      2 komik
      1 komiker
      3 komjölk
      1 komjölkallergi
      1 komjölksallergin
      1 komjölksproteinallergi
    153 komma
     18 kommande
      3 kommando
      1 kommenderade
      1 kommentar
      6 kommentarer
      1 kommentarerna
      1 kommentatorn
      3 kommenterade
      1 kommenterades
      4 kommenterar
    598 kommer
      1 kommersialisera
      1 kommersialiserade
      1 kommersialisering
      1 kommersialiseringen
      3 kommersiell
     10 kommersiella
      9 kommersiellt
      1 komminister
      1 kommissionär
      1 kommissionärerna
      9 kommissionen
      5 kommissionens
      1 kommisskläde
     82 kommit
      3 kommitté
      6 kommittén
     22 kommun
      8 kommunal
      7 kommunala
      1 kommunaliserades
      3 kommunalt
     16 kommunen
      1 kommunens
     13 kommuner
      4 kommunerna
      3 kommunernas
      1 kommuners
     12 kommunicera
      1 kommunicerande
      6 kommunicerar
     26 kommunikation
      4 kommunikationen
      1 kommunikationer
      1 kommunikationmetod
      8 kommunikationsavstånd
      2 kommunikationsavståndet
      1 kommunikationskontor
      1 kommunikationsleden
      3 kommunikationsproblem
      3 kommunikationssätt
      1 kommunikationsstörningar
      1 kommunikationssymtom
      1 kommunikationssystem
      1 kommunikationsteknologi
      1 kommunikationsteori
      1 kommunikationsunderlättande
      1 kommunikationsutrustning
      1 kommunikationsutrustningar
      2 kommunikativ
      1 kommunikativa
      2 kommunikativt
      2 kommuninvånarna
      1 kommuns
      1 kommutatorn
      1 komna
     12 komodo
      1 komodoensis
     11 komodovaran
     43 komodovaranen
      9 komodovaranens
     24 komodovaraner
      3 komodovaranerna
      1 komodovaranhona
      1 komorbid
      1 komorbida
      9 komorbiditet
      2 kompakt
      1 kompaktkassetten
      1 kompaniet
      1 kompaniets
      1 kompanisiffra
      1 kompanjon
      1 kompartementet
      1 kompartment
      2 kompartmentet
      4 kompartmentsyndrom
      1 kompartmentsyndromen
      1 kompatibelt
      3 kompatibilitet
      1 kompatibilitetsbedömningen
      1 kompatibla
      3 kompensation
      3 kompensationsmekanismer
      1 kompensatorisk
      9 kompensatoriska
      1 kompensatoriskt
     25 kompensera
      1 kompenserade
      4 kompenserar
      6 kompenseras
     13 kompetens
      1 kompetensbeviset
      1 kompetenscentrum
      2 kompetensen
      1 kompetenskrav
      2 kompetensutveckling
      2 kompetent
     28 komplement
      1 komplementaktivering
      2 komplementär
      1 komplementärmedicin
      1 komplementärmedicinsk
      1 komplementbrist
      1 komplementsystemet
      8 komplett
      4 kompletta
      8 komplettera
      1 kompletterad
      1 kompletterades
     13 kompletterande
      5 kompletterar
     12 kompletteras
      1 kompletterat
      2 komplettering
     31 komplex
     17 komplexa
      1 komplexet
      1 komplexitet
      4 komplexiteten
      9 komplext
      7 komplicerad
     13 komplicerade
      2 komplicerande
      2 komplicerar
      5 kompliceras
      6 komplicerat
     19 komplikation
      6 komplikationen
    109 komplikationer
      7 komplikationerna
      1 komplikationsfri
      1 komplikationsrisker
     15 komponent
      8 komponenten
     21 komponenter
      2 komponenterna
      2 komposit
      1 kompositer
      2 komposition
      1 kompositionen
      1 kompositioner
      1 kompositmaterial
      1 kompositörer
      1 komposteras
      5 kompresser
      5 kompression
      2 kompressioner
      1 kompressionerna
      4 kompressionsbehandling
      1 kompressionsstrumpor
      1 kompressorer
      7 komprimera
      2 komprimerad
      3 komprimerar
      9 komprimeras
      1 komprimerbara
      1 komprimering
      1 komprimeringsstället
      2 kompulsioner
      2 kompulsiva
      1 komvux
      1 kon
     56 kön
      1 konamikoden
      3 konästesier
      1 koncentrat
     32 koncentration
     35 koncentrationen
     24 koncentrationer
      3 koncentrationerna
      2 koncentrations
      3 koncentrationsförmåga
      1 koncentrationsförmågan
      1 koncentrationsgradiens
      2 koncentrationsgradient
      3 koncentrationsläger
      2 koncentrationslägren
      1 koncentrationsproblem
      1 koncentrationsprocess
      2 koncentrationsskillnaden
     17 koncentrationssvårigheter
      5 koncentrera
     22 koncentrerad
      7 koncentrerade
      4 koncentrerar
      5 koncentreras
      5 koncentrerat
      7 konceptet
      1 konception
      1 konceptualiseras
      1 koncernen
      1 koncernens
      1 koncis
      2 kondensationsreaktion
      1 kondensatorer
      4 kondenserar
      4 kondenseras
      1 kondenstorkskåp
      3 kondenstumlare
      8 kondition
      2 konditionen
      1 konditions
      1 konditionsidrott
      1 konditionskrävande
      1 konditionsträning
      1 konditorivaror
      1 kondoleanser
      1 kondolera
     23 kondom
      1 kondomanvändning
      1 kondomanvändningen
      9 kondomen
     16 kondomer
      1 kondomers
      1 kondomholkar
      1 kondrocyter
      1 kondrocyternas
      1 kondrodysplasi
      1 kondrodystropi
      6 kondrosarkom
      1 konduktionsafasi
     14 kondylom
     31 könen
      2 könens
      1 koner
      1 könet
      1 konferens
      1 konferensen
      1 konferenser
      3 konfessionella
      1 konfidensgrad
      2 konfidensintervall
      1 konfident
      1 konfiguration
      1 konfigurationsisomeren
      1 konfigurationsisomerer
      1 konfigureras
      1 konfirmation
      1 konfirmera
      1 konfirmerar
      1 konfiskera
     17 konflikt
      3 konflikten
     18 konflikter
      1 konfliktfritt
      1 konflikthypotesen
      3 konfliktlösning
      1 konfliktsituation
      1 konfokalmikroskopi
      1 konformade
      1 konformation
      1 konformationsändring
      2 konformationsförändring
      1 konformationsstress
      1 konformig
      1 konfrontativ
      2 konfrontativa
      1 konfucianska
      6 konfusion
      1 konfusionella
      1 konfusionen
      1 konfusionmedvetandesänkning
      2 kong
      4 kongenital
      1 kongenitala
      5 kongenitalt
      7 kongo
      5 kongokinshasa
      1 kongress
      1 kongressen
      1 kongresser
      1 kongressförhör
      1 konidieavsöndringen
      1 konidiebärare
      1 konidier
      2 konidierna
      2 koninklijke
      1 koniotomi
      3 konisk
      3 konjugation
      1 konjugera
      1 konjugerade
      1 konjugerar
      1 konjunktiv
      2 konjunktiva
      1 konjunktivit
      1 konkav
      1 konkava
      1 konkordansen
      1 konkordanta
      4 konkrement
     11 konkret
      7 konkreta
      1 konkretisera
      1 konkretiseras
      1 konkretisering
      1 konkubin
      1 konkurerade
      4 konkurrensen
      1 konkurrenskraft
      1 konkurrensutsatt
      2 konkurrent
      1 konkurrenter
      3 konkurrera
      6 konkurrerande
      3 konkurrerar
      1 konkurreras
      1 konkurrerat
      2 konkurs
      1 konkurser
      1 könlig
      1 könliga
      1 könligt
      2 könlös
      1 könlösa
      1 könlöst
      3 konnektivitet
      1 konnektiviteten
      1 könorganen
      1 konorski
      1 kons
      2 köns
      1 könsbehåring
      1 könsberoende
      1 könsbestämmande
      1 könsbunden
      1 könscell
      1 könscellen
     12 könsceller
      3 könscellerna
      1 könsdelar
      4 könsdelarna
      1 könsdifferentiering
      1 könsdifferentieringen
      1 könsdimorfism
      3 könsdrift
      1 könsdriften
      1 könsegenskaperna
     21 konsekvens
      6 konsekvensen
     34 konsekvenser
     11 konsekvenserna
      4 konsekvent
      1 konsekventa
     10 konsensus
      1 konsert
      2 konserter
      1 konserthus
      1 konserv
      1 konservatism
      6 konservativ
      5 konservativa
      1 konservative
      1 konservativt
      1 konservatorer
      1 konservburk
      1 konserven
      5 konserver
      3 konserverad
      1 konserveras
      2 konservering
      1 konserveringen
     15 konserveringsmedel
      1 könsfördelning
      2 könsfördelningen
      1 könshår
      1 könshormon
      6 könshormonbindande
     29 könshormoner
      7 könshormonerna
      1 könshormoners
      4 könsidentitet
      4 könsidentitetsstörning
      4 könsidentitetsstörningar
     11 konsistens
      3 konsistensen
      1 konsistensmedel
      1 konsistensökad
      1 könskaraktär
      6 könskarakteristika
      2 könskorrigerande
      3 könskorrigering
      1 könskörtel
      7 könskörtlar
      8 könskörtlarna
      1 könskromosmerna
      3 könskromosom
      1 könskromosomen
      5 könskromosomer
      2 könskromosomerna
      1 könskromosomparet
      1 könslig
      1 könsliga
      3 könsmogen
      6 könsmogna
      1 könsmognad
      2 könsmognaden
      1 könsmottagning
      1 könsneutral
      1 könsneutralt
      1 konsoliderades
      1 konsoliderar
      2 konsonant
      2 konsonanter
      1 konsonantföljder
     21 könsorgan
     16 könsorganen
      3 könsorganens
      2 könsorganet
      1 könsorgannjureörasyndrom
      1 konsortiet
      1 konsortium
      3 konspirationsteorier
      1 könsroller
      3 könssjukdom
      6 könssjukdomar
      2 könssjukdomarna
      2 könssjukdomen
      1 könsskiljande
      8 könsskillnader
      1 könsskillnaderna
      1 könsspecifik
      1 könsstörning
      1 könssträngstumörer
     12 konst
     31 konstant
      2 konstantinopel
     11 konstatera
      1 konstaterad
     13 konstaterade
      5 konstaterades
      1 konstaterandet
      6 konstaterar
      7 konstateras
      9 konstaterat
      9 konstaterats
      1 konstbefruktning
      1 konstellationer
      9 konsten
      1 konstfärdighet
      1 konstfibrer
      1 konstförståndiga
     16 konstgjord
      3 konstgjorda
      3 konstgjort
      1 konsthantverk
      2 konsthistoria
      2 konstig
      1 konstiga
      2 konstigt
      1 könstillhörighetslagen
      1 konstistensen
      4 konstitution
      1 konstitutionella
      1 konstitutiv
      1 konstlad
      5 konstnären
      7 konstnärer
      1 konstnärinnan
      4 konstnärliga
      3 konstnärligt
      1 konstnärskretsar
      1 konstnärskvarter
      1 konstnärssjäl
      1 konstnärssjälar
      1 konstrika
      4 konstruera
      1 konstruerad
      6 konstruerade
      6 konstruerades
      1 konstruerande
      2 konstrueras
      5 konstruerat
      6 konstruktion
      1 konstruktionell
      4 konstruktionen
      6 konstruktioner
      1 konstruktionsprincip
      1 konstruktionsprinciper
      4 konstruktiv
      2 konstruktivt
      1 konstruktören
      3 konstverk
      1 konstverken
      3 konstverket
      1 konsulent
      1 konsultarbete
      1 konsultation
      1 konsulter
      1 konsultera
      1 konsultfirma
      1 konsultverksamhet
      3 konsumenten
      9 konsumenter
      1 konsumentföreningen
      1 konsumentförpackning
      1 konsumentfrågor
      1 konsumentombudsmannen
      1 konsumentorganisationer
      1 konsumentpolitik
      2 konsumentprodukter
      1 konsumentrapporteringen
      4 konsumera
      1 konsumerade
     10 konsumerar
      3 konsumeras
      2 konsumerat
      2 konsumerats
      1 konsumering
      1 könsumgänge
      1 konsumism
     27 konsumtion
      4 konsumtionen
      1 konsumtionsfaser
      1 konsumtionsvaror
      2 könsutveckling
      1 könsutvecklingen
    174 kontakt
     18 kontakta
      1 kontaktade
      2 kontaktallergener
     12 kontaktallergi
      1 kontaktallergin
      1 kontaktallergiskt
     10 kontaktas
      1 kontaktaureoler
      1 kontaktbehandling
      2 kontaktdermatit
      6 kontakteksem
      6 kontakten
      9 kontakter
      1 kontaktgoniometern
      2 kontaktlins
      1 kontaktlinsen
     12 kontaktlinser
      2 kontaktlinserna
      1 kontaktlinsvätskor
      1 kontaktmetamorfos
      1 kontaktperson
      1 kontaktpunkten
      1 kontaktsmitta
      2 kontaktspårning
      1 kontaktstörning
      1 kontakttid
      1 kontaktyta
      1 kontaktytor
      6 kontamination
      1 kontaminationsfrekvensen
      2 kontaminerad
      3 kontaminerade
      1 kontaminerar
      1 kontamineras
      1 kontaminerat
      2 kontemplation
      2 kontemplationen
      1 kontemplativa
      3 kontext
      1 kontinens
      1 kontinent
      3 kontinenten
      4 kontinenter
      1 kontinenterna
     10 kontinuerlig
      3 kontinuerliga
     32 kontinuerligt
      2 kontinuitet
      1 kontinuumet
      2 kontoinnehavare
      1 kontoinnehavaren
      1 kontoinnehavarens
      1 konton
      4 kontor
      1 kontorsanställda
      1 kontorsmaskin
      1 kontorsmiljö
      1 kontorspersonal
      1 kontorsrum
      3 kontot
      2 kontra
      1 kontrafobier
      5 kontrahera
      6 kontraherar
      1 kontraherardras
      1 kontrahering
      1 kontraindicerad
      1 kontraindikation
      1 kontraindikationer
      7 kontrakt
      5 kontraktet
      1 kontraktil
      8 kontraktion
      3 kontraktionen
      2 kontraktioner
      1 kontraktsmålet
      1 kontraktsslut
      1 kontraktuell
      1 kontrakturer
      5 kontralateral
      1 kontralaterala
      5 kontrast
      2 kontrasten
      1 kontraster
      1 kontrastförluster
      8 kontrastmedel
      3 kontrastmedlet
      2 kontraströntgen
      1 kontrastskillnad
      3 kontrastvätska
      1 kontratenorer
      1 kontraterrorism
      1 kontraterroriststyrkor
     93 kontroll
      1 kontrollåtgärder
      9 kontrollen
     13 kontroller
     45 kontrollera
     17 kontrollerad
     15 kontrollerade
      1 kontrollerades
     21 kontrollerar
     22 kontrolleras
      3 kontrollerat
      4 kontrollerna
      2 kontrollgrupp
      2 kontrollgruppen
      3 kontrollgrupper
      2 kontrollmekanism
      1 kontrollmekanismer
      1 kontrollodla
      1 kontrollorgan
      1 kontrollsummor
      1 kontrollverksamhet
      6 kontrovers
      2 kontroversen
      4 kontroverser
     15 kontroversiell
      5 kontroversiella
     14 kontroversiellt
      1 kontur
      3 konturer
      1 konung
      2 konvalescens
      1 konvalescentsera
      1 konvaljväxter
      1 konvektion
      1 konvent
     16 konvention
      8 konventionell
      9 konventionella
     20 konventionen
      1 konventioner
      2 konventionerna
      1 konversation
      2 konversationell
      2 konversationen
      5 konvertera
      1 konverterades
      1 konverterar
      1 konverteras
      1 konvertering
      1 konverteringen
      1 konvex
      2 konvexa
      3 konvulsioner
      1 konvulsiv
      1 konvulsiva
      1 konvulsivisk
     15 konzo
      1 konzoutbrott
      1 kooperativ
      3 koordination
      1 koordinationen
      1 koordinationsförmågan
      4 koordinera
      1 koordinerad
      1 koordineras
      2 koordinerat
      4 köp
     28 köpa
      1 köpande
      1 köpare
      2 köparen
      1 köparna
      7 köpas
      1 köpcentret
      1 köpekontraktet
      5 köpenhamn
      1 köpenhamns
      5 köper
      1 köpet
      6 kopia
      2 kopiera
      1 kopierade
      1 kopierar
      1 kopieras
      1 köping
      4 kopior
      1 kopiorna
      1 kopolymer
      2 kopp
      1 koppa
     21 koppar
      1 kopparacetat
      1 kopparbaserat
     11 kopparbrist
      1 kopparcyanid
      1 kopparhaltigt
      5 kopparhuvud
      2 kopparintag
      1 kopparmolekyler
      1 kopparn
      2 kopparnivåerna
      1 kopparns
      1 kopparoxid
      1 kopparplåtar
      1 koppärr
      4 kopparspiral
      1 kopparspiraler
      1 kopparstenåldern
      1 koppartransporterande
      1 kopparyxa
      1 koppas
      1 koppeltvång
     11 koppen
      1 kopphorn
      6 koppla
     13 kopplad
     27 kopplade
      1 kopplades
      6 kopplar
     29 kopplas
     21 kopplat
      4 kopplats
     38 koppling
      8 kopplingar
      2 kopplingarna
     19 kopplingen
      1 kopplingsarbete
      1 kopplingspunkt
      1 kopplingspunkten
      1 kopplingspunkter
      1 kopplingsstation
      7 koppning
      1 koppor
      1 kopporna
      1 kopra
      5 koprolali
      1 koproporfyrinogen
      1 kopropraxia
      1 kopros
      1 koprostas
      2 köps
      1 köpt
      4 köpte
      3 köptes
      1 kopulation
      1 kopulationen
      1 kopulera
     17 kor
     10 kör
     17 köra
      1 korall
      2 korallbär
      1 korallbuskar
      1 korallbusksläktet
      3 koralldjur
      1 korallrev
      5 koranen
      1 [koranen
      2 köras
      1 körbana
      1 körbanan
      1 körbeteende
      1 korda
      1 kördugligheten
      7 korea
      1 koreahalvön
      1 koreakriget
      1 koreansk
      1 koreanska
      1 koreografi
      1 körfältsförändringar
      1 korg
      2 korgarna
      2 korgblommiga
      1 körhandtagen
      1 koriander
      1 koriomeningitisvirus
      1 korionbiopsi
      1 koriongonadotropin
      1 koriskt
      2 körkort
      1 korkskruv
      1 körlar
      3 korm
      1 kormen
      1 kormfluga
      1 kormflugans
     12 korn
      1 kornea
      1 kornealmikroskop
      1 kornealreflexen
      1 kornen
      1 kornets
      1 korniga
      1 kornigt
      2 körning
      1 körnskörtlarna
      1 koronarangiografi
      1 koronarkärlssjuka
      1 koronarstentar
      1 koronartrombos
      1 koronis
      1 korpavföring
      2 korpulens
      1 korregeras
     33 korrekt
     11 korrekta
      2 korrektion
      3 korrektionsglas
     14 korrelation
      3 korrelationen
      1 korrelationer
      2 korrelationsanalyser
      6 korrelera
      1 korrelerad
      2 korrelerade
     21 korrelerar
      1 korrelerat
      1 korrellerar
      1 korrespondens
      1 korresponderande
      1 korresponderar
     13 korrigera
      1 korrigerad
      1 korrigerade
      2 korrigerande
      3 korrigerar
      6 korrigeras
      1 korrigerat
      1 korrigerats
      5 korrigering
      1 korrigeringsalternativet
      1 korrodering
      1 korrosion
      1 korrosionens
      1 korrosivt
      1 korrossion
      1 korrupta
      1 korruption
      3 kors
      2 körs
      3 korsa
      1 korsade
      7 korsallergi
      4 korsande
      7 korsar
      2 korsas
      1 korsat
      1 körsbärskärnor
      2 körsbärsliknande
      1 körsbärsstora
      1 körsbärstomater
      1 korsbinds
      3 korsblommiga
      1 korsbunden
      1 korsdrag
      1 korselett
      1 korseletten
      1 korseletter
      2 korset
     13 korsett
      1 korsettanvändandet
     24 korsetten
      2 korsettens
     14 korsetter
      1 korsettering
      1 korsetteringen
      2 korsetterna
      1 korsettindustrin
      1 korsettliknande
      2 korsettliv
      1 korsettlivet
      1 korsettmodet
      1 korsettyper
      1 korsfäst
      4 korsika
      1 korslagda
      1 korslänkas
      3 korsning
      2 korsningar
      4 korsningen
      1 korspollinering
      1 korsreagerande
      1 korsreagerar
      1 korsreaktion
      1 korsreaktioner
      1 korsreaktiva
      2 korsryggen
      2 korståg
      1 korstestat
      1 korstolerant
      1 korsväg
     94 kort
     42 korta
      1 kortänden
      2 kortar
     60 kortare
      1 kortast
      2 kortaste
      9 körtel
      1 körtelcancer
      2 körtelcell
      1 körtelceller
      1 körtelcellerna
      6 körtelfeber
      3 körtelgångar
      6 körteln
      1 körtelpaket
      1 körtelparti
      1 körtelsvulst
      1 körteltäta
      2 körtelvävnad
      4 körtelvävnaden
      1 körtelvävnaderna
      1 korten
      1 kortex
      1 kortfattade
      2 korthet
      1 korthuvud
      2 kortikal
      4 kortikala
      2 kortikosteroid
     14 kortikosteroider
      3 kortikotropin
      2 kortikotropinfrisättande
     26 kortisol
      1 kortisoldehydroepiandrosteronkvoten
      1 kortisoler
      1 kortisolinjektion
      1 kortisolnivån
      1 kortisolutsöndring
      1 kortisolvärdena
     23 kortison
      3 kortisonbehandling
      1 kortisonet
      1 kortisonhaltiga
      2 kortisoninjektioner
      1 kortisonkräm
      2 kortisonpreparat
      2 kortisonsalva
      1 kortisonsalvor
      2 kortisontabletter
      1 kortkedjiga
     32 körtlar
     11 körtlarna
      2 körtlarnas
      1 körtlarutsöndringsmekanismer
      1 körtlens
      1 kortlivad
      3 kortlivade
      1 kortroman
      1 körts
      1 kortsiktig
      3 kortsiktiga
      4 kortsiktigt
      1 kortsiktligt
      1 kortskalle
      1 kortslutningar
      2 kortspel
      2 korttidsanvändning
      1 korttidsbehandling
      1 korttidsfasta
      1 korttidsförvara
      2 korttidsminne
      1 korttidsterapi
     15 kortvarig
      6 kortvariga
     10 kortvarigt
      1 kortväxthet
      2 kortverkande
      1 kortvuxenhet
      3 korv
      1 korvskinn
      2 kos
      2 kosher
      1 kosherkrav
      5 kosjukan
     10 kosmetika
      2 kosmetikaföretag
      1 kosmetikatester
      1 kosmetikavärlden
      1 kosmetikdirektivet
      1 kosmetiktillverkare
      7 kosmetisk
     21 kosmetiska
      5 kosmetiskt
      1 kosmiska
      1 kosmologi
      1 kosmologiskt
      4 kosmos
     91 kost
      3 kosta
     11 kostar
      2 kostat
      2 kostbehandling
      1 kostbehandlingen
      1 kostbeteende
      1 kostbyte
      2 kostcirkeln
      1 kostcirkelns
     26 kosten
      4 kostens
      2 kostfaktorer
      2 kostfiber
      1 kostfibrer
      1 kostförändring
      1 kosthålling
     22 kosthållning
      2 kosthållningen
      1 kosthälsoinformation
      1 kostinformation
      1 kostinnehåll
      1 kostintag
      1 kostintaget
      1 kostkorrigeringar
     12 kostnad
     13 kostnaden
     20 kostnader
      5 kostnaderna
      1 kostnadseffektanalys
      2 kostnadseffektiv
      2 kostnadseffektiva
      1 kostnadseffektivare
      4 kostnadseffektivt
      2 kostnadsfri
      1 kostnadsfria
      3 kostnadsfritt
      1 kostodiafragmala
      1 kostomläggning
      1 kostplanen
      1 kostprogram
      4 kostråd
      1 kostråden
      2 kostrådgivning
      1 kostreglering
      1 kostrekommendationer
      1 kostrekommendationerna
      2 kostrelaterade
      5 kostsam
      1 kostsamma
      1 kostsamt
     11 kosttillskott
      3 kostvanor
      1 kostverk
      2 kostym
      1 kostymgalge
      1 kotan
      1 kotknackare
      1 kotkompression
      7 kotodama
      5 kotor
      6 kotorna
      4 kototama
      1 kototamans
      1 kotpelare
      1 kotpelaren
      1 kotsegment
     52 kött
      1 köttäggmejeriprodukter
      1 kottarna
      4 köttätande
      1 köttätandet
      1 köttätare
      1 köttberget
      1 köttbiten
      1 kotte
      1 kottepalmer
     10 köttet
      1 köttfärs
      3 köttig
      5 köttiga
      3 köttklister
      1 köttklöven
      2 köttprodukter
      1 köttprov
      1 köttsaften
      2 köttstycken
      1 kousha
      1 kousis
      1 kovalenta
      1 kövarning
      5 kpa
      1 kpenumoniae
      7 kpneumoniae
     18 kr
      2 krabba
      1 krabbakräfta
      2 kraepelin
      1 kraepelins
      1 krafftebing
     44 kraft
      2 kräfta
      1 kraftdjur
      1 kräftdjur
      7 kraften
     12 krafter
      5 krafterna
      1 kraftfältet
      1 kraftfoder
      5 kraftfull
      4 kraftfulla
      1 kraftfullare
      1 kraftfullaste
      3 kraftfullt
     82 kraftig
     48 kraftiga
     14 kraftigare
      1 kraftigast
      3 kraftigaste
    132 kraftigt
      2 kraftledningar
      1 kraftlös
      4 kraftlöshet
      1 kraftnedsättning
      1 kraftpåverkningar
      1 kraftproducerande
      1 kraftprov
      1 kräftriket
      1 kraftstärkande
      1 kraftuttryck
      1 kraftvektorn
      1 kraftverkan
      1 kragen
     10 kräkas
      2 kraken
      1 kräkformen
      1 kräkmedlen
     24 kräkning
     73 kräkningar
      1 kräknötsväxter
      4 kräkreflexen
      1 kräkreflexer
      5 kräks
      1 kräktoxinet
      1 kräkts
      4 kräldjur
     10 kräm
      1 kramades
      1 kramas
      1 krämen
      8 krämer
      1 krämfärgat
      1 kramning
     10 kramp
      2 krämpa
      2 krampaktig
     16 krampanfall
      1 krampartad
      1 krampbenägenhet
      1 krampbenäget
      1 krampen
     30 kramper
      3 kramperna
      1 krampkänslor
      2 kramplösande
      1 krämpor
      1 krampspasmlösande
      1 kramptillstånd
      1 krånglande
      2 krångliga
      1 krängning
      1 kranialnerv
      1 kranialnerven
      2 kranialnerver
      3 kranialnerverna
      1 kraniekapaciteter
      1 kraniella
      4 kranier
     10 kraniet
      1 kräningar
      3 kraniofaryngiom
      1 kranium
      1 kränka
      1 kränkande
      1 kränker
      2 kränkning
      1 kränkt
      5 krans
      2 kransar
      1 kransbindning
     15 kranskärl
      3 kranskärlen
      2 kranskärlet
      1 kranskärlsoperationer
      4 kranskärlsröntgen
      1 kranskärlssjukdom
      1 kranvatten
      1 kräppat
      1 kras
      1 krasis
      1 kräsna
      1 krater
     84 krav
      1 kräv
     15 kräva
      1 kravallbekämpning
      1 kravallsköldar
      7 krävande
     10 krävas
      9 krävde
      8 krävdes
     23 kraven
    144 kräver
      8 kravet
      2 kravitz
      1 kravmärkt
      1 kravnivå
    183 krävs
      2 krävt
      1 krazy
      1 kreatin
      2 kreatinin
      1 kreatininstegring
      4 kreatinkinas
      1 kreativ
      2 kreativa
      3 kreativitet
      2 kreativiteten
      1 kreatur
      1 kreaturskötseln
      1 kreditbanken
      1 kreditinstitut
      1 krematorienbauers
      1 krematorier
      1 kremerades
      1 kremlor
      1 krenitism
      1 kreosot
      5 kresol
      1 kresolens
      2 kreta
      4 kretek
      3 kretin
      6 kretinism
      2 krets
      1 kretsa
      1 kretsade
     13 kretsar
      4 kretsen
      5 kretslopp
     11 kretsloppet
      1 kretsloppstänkande
      1 kretzschmaria
     15 krig
      1 krigarkulturer
      1 krigen
      7 kriget
      1 krigförande
      3 krigföring
      1 krigsbrott
      1 krigsbyten
      2 krigsdimma
      2 krigsfångar
      1 krigsförbrytelse
      1 krigsguden
      1 krigsinvalider
      1 krigskirurg
      1 krigsmakten
      1 krigsneuros
      1 krigsproduktion
      1 krigståg
      1 krigsveteraner
      2 krigszoner
      1 krikofaryngeusmuskeln
      4 krim
      1 kriminalfilmer
      2 kriminaliserade
      1 kriminaliserades
      1 kriminaliserar
      1 kriminaliserat
      1 kriminalisering
      1 kriminaliseringen
      6 kriminalitet
      1 kriminalpoliser
      2 kriminalvården
      3 kriminell
     13 kriminella
      1 kriminellas
      1 kriminelle
      4 kriminellt
      1 kriminologen
      1 kriminologi
      1 kriminologisk
    175 kring
      1 kringfarande
      1 kringgår
      4 kringliggande
      1 kringresande
      2 kringströdda
      1 krinolin
      6 kris
      2 krisberedskap
      1 krisen
      7 kriser
      1 krisfyllda
      1 krishantering
      1 krishnamacharya
      1 krisreaktioner
      1 krissituationer
      1 krisstöd
      3 kristall
      1 kristallation
      2 kristallbildningen
      1 kristallblad
      5 kristallen
     23 kristaller
      2 kristallerna
      1 kristallernas
      1 kristallfasens
      2 kristallin
      2 kristallina
      2 kristallinskt
      1 kristallint
      1 kristallisation
      2 kristalliserad
      2 kristalliserade
      2 kristalliserar
      1 kristalliseras
      2 kristalliserat
      1 kristalliter
      1 kristallmassa
      1 kristallografin
      1 kristallpulver
      1 kristallscintillatorer
      1 kristallsjukan
      6 kristallstruktur
      6 kristallsystem
      1 kristallytan
      1 kristallytor
      1 kristallytorna
      2 kristallytornas
      8 kristen
      4 kristendom
      7 kristendomen
      4 kristendomens
      1 kristendomskritik
      1 kristian
      1 kristianstad
      1 kristider
      2 kristina
     25 kristna
      1 kristofer
      9 kristus
      2 krita
     31 kriterier
     14 kriterierna
      4 kriteriet
      4 kriterium
      1 kritierium
     52 kritik
      1 kritikdebatt
     16 kritiken
     22 kritiker
     10 kritikerna
      1 kritisera
      5 kritiserade
      1 kritiserades
      3 kritiserar
      2 kritiseras
      2 kritiserat
     15 kritiserats
      9 kritisk
     14 kritiska
      5 kritiskt
      2 kritpipor
      1 kro
      2 krock
      2 krocka
      1 krockar
      2 kroenke
      2 krogar
      1 krogen
      2 krok
      6 krökar
      1 kröken
      4 kröker
      3 krokidolit
      3 krokiga
      7 krökning
      1 krökningen
      1 krökningens
      1 kroknosa
      1 krokodiler
      1 kröks
      3 krökt
      3 krökta
      1 krokusar
      1 krokusarna
      1 krokusliljesläktet
      5 krom
      1 kromallergi
      1 kromat
      1 kromatin
      1 kromatinet
      2 kromatinremodellering
      6 kromatografi
      1 kromatografin
      3 kromatografiska
      1 kromiiioxid
      1 kromkoboltlegering
      1 kromoglikat
     28 kromosom
      4 kromosomala
      2 kromosomalt
      3 kromosomavvikelse
      1 kromosomavvikelsen
      8 kromosomavvikelser
      1 kromosombild
      6 kromosomen
     19 kromosomer
      7 kromosomerna
      1 kromosomernas
      1 kromosomfel
      1 kromosomförändring
      1 kromosomförändringar
      5 kromosompar
      1 kromosomregioner
      1 kromosomrubbning
      1 kromosomrubbningssyndrom
      1 kromosomtal
      1 kromosomtypen
      1 kromosomuppsättning
      1 kromosomuppsättningar
      1 kromosomuppsättningen
      1 kromsalter
      1 kromsyra
      6 krona
      1 kronägg
      7 kronan
      1 kronans
      8 kronblad
      6 kronbladen
      1 kronbladslika
      1 kronbladsliknande
      1 kronchakrat
      1 kronebrott
      1 kronflikarna
      1 krönika
      2 kronisering
    135 kronisk
     46 kroniska
     17 kroniskt
      1 kronobergs
      1 kronologi
      1 kronologin
      2 kronologisk
      1 kronologiska
      1 kronologiskt
     25 kronor
      1 kronordag
      2 kronorsemblem
      2 kronoterapi
      2 kronotyp
      1 kronotypen
      1 kronstam
      1 kropdel
     79 kropp
     18 kroppar
      3 kropparna
      1 kroppars
    725 kroppen
    248 kroppens
      1 kroppentemperaturen
      1 kroppentumören
      1 kroppenupplevelser
      1 kroppfunktioner
      5 kropps
      1 kroppsaktivitet
      2 kroppsansträngning
      1 kroppsansträngningar
      1 kroppsarbetare
      1 kroppsarbete
      1 kroppsbehandling
      2 kroppsbehåring
      1 kroppsbelastning
      1 kroppsbild
      1 kroppsburet
      2 kroppsbyggnad
     18 kroppsdel
     34 kroppsdelar
      4 kroppsdelarna
     10 kroppsdelen
      1 kroppsdels
      2 kroppsegen
      2 kroppseget
      1 kroppsegment
      3 kroppsegna
     20 kroppsfett
      1 kroppsfetter
      1 kroppsfettet
      3 kroppsform
      3 kroppsformen
      3 kroppsfrämmande
      1 kroppsfunktion
      8 kroppsfunktioner
      1 kroppsgena
      3 kroppshålan
      1 kroppshålans
      1 kroppshåligheter
      3 kroppshållning
      1 kroppshålor
      1 kroppshålorna
      3 kroppshalva
      2 kroppshalvan
      1 kroppshår
      1 kroppsideal
      1 kroppsjuveler
      1 kroppskännedom
      1 kroppskännedomsövningar
      3 kroppskontakt
      1 kroppslägen
      2 kroppslängd
      1 kroppslängden
     26 kroppslig
     24 kroppsliga
      1 kroppsligkinestetisk
      5 kroppsligt
      6 kroppslukt
      4 kroppslukten
      2 kroppsmålning
      2 kroppsmassa
      1 kroppsmått
      1 kroppsmåtten
      1 kroppsmedvetenhet
      1 kroppsmodifikation
      1 kroppsöppning
      2 kroppsöppningar
      2 kroppsöppningarna
      1 kroppsorganens
      3 kroppsövningar
      1 kroppspiercingen
      1 kroppsposition
      1 kroppsproportioner
      2 kroppspsykoterapi
      6 kroppspulsådern
      1 kroppsrengöring
      1 kroppsrörelsen
      3 kroppsrörelser
      1 kroppssammansättning
      3 kroppssegment
      1 kroppsskador
      4 kroppsspråk
      2 kroppsställning
      1 kroppsställningar
      2 kroppsstorlek
      1 kroppssvettningar
      1 kroppssymmetrin
     31 kroppstemperatur
     18 kroppstemperaturen
      2 kroppstemperaturer
      1 kroppstempertur
      1 kroppsterapimetoder
      2 kroppstyp
      4 kroppsundersökning
      2 kroppsundersökningar
      5 kroppsuppfattning
      2 kroppsuppfattningen
      1 kroppsutsmyckning
      3 kroppsväggen
      5 kroppsvärme
      3 kroppsvätska
      1 kroppsvätskan
     12 kroppsvätskor
      6 kroppsvätskorna
      1 kroppsvätskornas
      1 kroppsvävander
      6 kroppsvävnad
      1 kroppsvävnaden
     18 kroppsvikt
      4 kroppsvikten
      1 kroppsvisitation
      1 kroppsyta
      2 kroppsytan
      1 kroppvätskor
      5 krossade
      1 krossar
      2 krossas
      3 krossat
      1 krosskador
      1 krosslink
      1 krosslinkade
      1 krosslinkare
      1 krotonolja
      1 krs
      1 krugerrand
      1 kruka
      1 krukan
      1 krukor
      6 krukväxt
      4 krukväxter
      1 krumtarm
      2 krumtarmen
      2 krupp
      1 krusbär
      1 krycka
      1 kryckan
      2 kryckor
      4 krydda
      1 kryddiga
      1 kryddmått
      3 kryddnejlika
      4 kryddor
      1 kryddörter
      1 kryddsill
      1 kryddsmak
      1 kryddstark
      1 krylovii
      4 krympa
      2 krymper
      1 krymplingar
      1 krympning
      4 kryonik
      1 kryoniker
      2 kryoteknik
      4 krypa
      7 krypande
      4 kryper
      2 krypningskänslor
      1 krypstadium
      1 kryptogamer
      1 kryptokockantigen
      5 kryptokockmeningit
      1 kryptor
      5 kryptorkism
      1 kryptorna
      1 kryptos
      2 kryptosporidios
      1 kryptozoologi
      7 krysotil
      1 kryssen
      1 kryssmärke
      1 kryssmärkena
      1 kryssmärket
      1 krysta
      1 krystar
      2 krystas
      1 krystning
      1 krystningar
      1 krystningsskedet
      1 krystningstiden
      1 krystvärkarna
      1 ksh
      1 kspecifika
      2 k�t
      1 kth
      1 ktha
      1 ktmtranssexuella
      3 kts
      2 kuba
      1 kubikmeter
      1 kubikmillimeter
      1 kubisk
      3 kubiska
      2 kubiskt
      3 kubmaneter
      1 kubtest
      1 kucinich
      6 kuddar
      2 kudde
      1 kuddformad
      4 kuff
      1 kuffas
      3 kuffen
      1 kuffvätskemängden
      1 kugler
      2 kula
      1 kulformade
      3 kull
      1 kullar
      1 kullstorleken
      7 kulmen
      1 kulminerade
      3 kulor
      1 kulör
      1 kulörer
      1 kulört
      2 kulörta
      1 kulsiltyperna
      1 kulspruta
      1 kulsprutepistol
      1 kulsprutor
      1 kult
      2 kultivarer
      1 kultiverade
      1 kultstatus
     24 kultur
      1 kulturarvet
      1 kulturberoende
      2 kulturbundna
      1 kulturcentra
      1 kulturchock
      4 kulturell
     21 kulturella
      5 kulturellt
     13 kulturen
      1 kulturens
     36 kulturer
      1 kulturerna
      1 kulturers
      2 kulturhistoria
      1 kulturjord
      1 kulturkrock
      1 kulturmedicin
      1 kulturnämnderna
      1 kulturref
      1 kulturrelaterad
      1 kultursektorn
      1 kultursfärerna
      2 kulturspecifika
      1 kulturspecifikt
      1 kulturväxt
      1 kulturväxter
      1 kulturvetenskap
      2 kumarin
      1 kumarintyp
      2 kumen
      1 kumenprocessen
      1 kumlingesjukan
      2 kumulativ
      1 kunaindianerna
      1 kund
      2 kunda
      1 kundali
     11 kundalini
      1 kundalinienergin
      1 kundalinigudinnan
      4 kundalinikraften
      1 kundalinisyndromet
      1 kundaliniterapi
      1 kundalinivaknande
      5 kundaliniyoga
      2 kundaliniyogan
      1 kundbasen
    255 kunde
      6 kunden
      1 kundens
      7 kunder
      1 kunderna
      1 kundernas
      2 kunders
      1 kundvänligare
     10 kung
      2 kungafamiljen
      1 kungahus
      2 kungahusen
      1 kungakrona
      1 kungakronor
      1 kungamakten
      1 kungar
      8 kungen
      1 kungens
      1 kungl
      1 kunglig
      5 kungliga
      1 kungligheter
      1 kungligt
      1 kungörelser
      2 kungsholmsloka
      1 kungskobra
      1 kungsörs
      1 kunkurrera
    433 kunna
     70 kunnat
      1 kunnig
      2 kunniga
     80 kunskap
     15 kunskapen
     21 kunskaper
      4 kunskaperna
      1 kunskaps
      1 kunskapsbas
      1 kunskapsdatabas
      1 kunskapsdisciplinerna
      2 kunskapsfält
      2 kunskapsinhämtning
      1 kunskapskrav
      1 kunskapsläget
      2 kunskapsnivå
      1 kunskapsområdena
      1 kunskapsområdet
      1 kunskapsöversikt
      1 kunskapsteori
      1 kunskapsunderlag
      2 kupa
      2 kupan
      1 kupbredden
      1 kupmått
      1 kupning
      2 kupor
      1 kuporna
      4 kupstorlek
      2 kupstorlekar
      2 kupstorleken
      6 kur
      1 kurativ
      4 kurator
      2 kuratorer
      1 kurbma
      1 kurbrandenburska
      1 kurdiska
      5 kuren
      2 kurer
      4 kurera
      1 kurerande
      1 kurerna
      1 kurett
      1 kurhmä
      2 kurhus
      1 kurhusavdelningar
      1 kurhusavgiften
      4 kuriosa
      1 kuriosakunskaper
      1 kuriositet
      5 kurkumin
      1 kurmetod
      1 kurort
      1 kurortens
      1 kurorter
      1 kurorterna
      1 kurrande
      5 kurs
      1 kursavgiften
      1 kursens
      4 kurser
      1 kurserna
      1 kursplan
      1 kursutbildning
      3 kurt
      1 kurtis
      1 kurtiseringsuppgörelser
      1 kuru
      6 kurva
      5 kurvan
      1 kurvform
      1 kurvig
      3 kurvor
      1 kurvorna
      1 kurze
      1 kushi
      1 kusin
      1 kusinäktenskap
      1 kusinerna
      1 kusingifte
      1 kusingiften
      1 kuske
      1 kuskohygrin
      1 kussmauls
      2 kust
      1 kustbefolkningen
      1 kusten
      2 kuster
      1 küster
      1 kusterna
      1 kustlandskap
      1 kustlinje
      1 kustmarkens
      1 kustområden
      1 kustområdet
      1 kustsediment
      2 kusttrakter
      1 kustvatten
      1 kutan
      2 kutluk
      1 kuusisito
      1 kuusisto
      1 kuvalayananda
      1 kuvert
      3 kuvös
      4 kuvösen
      3 kuvöser
      1 kuvöserna
      1 kuvösvården
      1 kuwait
      3 kv
      1 kvacka
      5 kvacksalvare
      8 kvacksalveri
      1 kvacksalveribehandlingar
      3 kvacksalverilagen
      1 kvaddlar
      2 kvadrat
      1 kvadratisk
      1 kvadratkilometer
      2 kvadratmeter
      1 kvadrivalent
      1 kval
      1 kvalificera
      7 kvalificerad
      3 kvalificerade
      2 kvalificerar
      3 kvalificerat
      2 kvalitativ
      1 kvalitativa
      2 kvalité
      4 kvalitén
     23 kvalitet
      7 kvaliteten
      3 kvaliteter
      1 kvalitetsbedömning
      1 kvalitetsfaktor
      2 kvalitetsfaktorn
      1 kvalitetshöjning
      1 kvalitetsindikationer
      1 kvalitetsindikator
      2 kvalitetsjusterade
      1 kvalitetskontrollen
      1 kvalitetskrav
      1 kvalitetskriterierna
      1 kvalitetsmärkning
      1 kvalitetsmärkt
      1 kvalitetsnivå
      1 kvalitetsproblem
      1 kvalitetssäkring
      1 kvalitetssäkringskrav
      1 kvalitetssegment
      1 kvalitetssynpunkt
      4 kväll
      1 kvällar
      2 kvällarna
      7 kvällen
      1 kvällstid
      6 kvalster
      3 kvalsterburna
      1 kvantal
      1 kvantifieras
      1 kvantifierbara
      2 kvantifiering
      4 kvantitativ
      1 kvantitativt
      3 kvantitet
      2 kvantiteten
      3 kvantiteter
      1 kvantitetsbetyg
    133 kvar
      1 kvarblir
      2 kvardröjande
      1 kvardröjd
      2 kvardröjer
      2 kvarhållande
      2 kvarhållas
      1 kvarhållning
      1 kvarhöll
      1 kvarka
      1 kvarkatetrar
      1 kvarlämnade
      1 kvarlämnas
      5 kvarleva
      5 kvarlevor
      1 kvarlevorna
      8 kvarliggande
     11 kvarstå
      6 kvarstående
     21 kvarstår
      2 kvarstod
      1 kvart
      2 kvartalet
      1 kvartalslinser
      2 kvartär
      1 kvarteret
      1 kvarts
      1 kvartskristall
      1 kvartspartiklarna
     11 kvarvarande
      1 kvasibiologi
      1 kvastklassifikation
      1 kvastlika
      1 kvatemberveckorna
      2 kväva
      2 kvävande
      1 kvävas
      1 kvävda
     16 kväve
      1 kväveavskiljningen
      1 kvävebas
      1 kvävebasen
      2 kvävedioxid
      1 kvävehalt
      1 kvävehaltig
      1 kvävehaltiga
      1 kvävehaltigt
      1 kväven
      3 kvävenarkos
      1 kvävenärsalter
      8 kväveoxid
      1 kväveoxidul
      1 kväver
      2 kväverik
      1 kvävet
      1 kvävetrijodid
      1 kvävetrijodidkristaller
      1 kväveupptaget
      6 kvävgas
      1 kvävgasen
     12 kvävning
      1 kvävningskänslor
      1 kvesved
      1 kvicka
      1 kvicknar
      2 kvickrot
     26 kvicksilver
      1 kvicksilverånga
      2 kvicksilverförgiftning
      1 kvicksilverhalt
      1 kvicksilveroxid
      1 kvicksilversalva
      1 kvicksilversalvor
      1 kvicksilvertekniken
      1 kvicksilvertermometrar
      3 kvicksilverutsläpp
      1 kvicksilvret
      1 kvickt
     87 kvinna
      1 kvinnaman
    155 kvinnan
      1 kvinnanflickan
     66 kvinnans
      9 kvinnas
      2 kvinnatillman
     17 kvinnlig
     47 kvinnliga
      1 kvinnlighet
      8 kvinnligt
      1 kvinno
      7 kvinnobröst
      1 kvinnobrösten
      1 kvinnodräkten
      1 kvinnofientligt
      1 kvinnoförtryck
      1 kvinnohänder
      1 kvinnoklinik
      2 kvinnokliniker
      1 kvinnokropp
    580 kvinnor
      1 kvinnorättsorganisation
     26 kvinnorna
      2 kvinnornas
      1 kvinnoröster
     26 kvinnors
      1 kvinnosjukvård
      1 kvinnosynen
      1 kvinnoyrke
      1 kvint
      1 kvisslor
      2 kvist
      2 kvistar
      1 kvistarna
      2 kvisten
      5 kvitamin
      2 kvitt
      1 kvittblivningsvolymen
      1 kvitten
      7 kvot
      1 kvotberäkning
     10 kvoten
      2 kvoter
      1 kwakiutul
      1 kwanghung
      1 kwangoområdet
      4 kwashiorkor
      1 kyanol
      1 kyasanur
      9 kyckling
      1 kycklingar
      1 kycklingbröst
      1 kycklingskinn
      1 kycklingsoppa
     28 kyla
      1 kylan
      2 kylande
      8 kylarvätska
      1 kylbox
      1 kylen
      3 kyler
      1 kylförvaras
      1 kylig
      1 kyliga
      5 kyligt
      1 kylklampar
      3 kylmedel
      1 kylmekanism
      6 kylning
      1 kylomikroner
      1 kylös
      1 kylpåse
      1 kylpåsen
      1 kylrum
      1 kyls
      5 kylskåp
      1 kylskåpkylrum
      1 kyltorn
      1 kylus
      1 kylvaror
      1 kylväska
      4 kylväskan
      2 kylväskor
      2 kylväskorna
      1 kymotrypsinogen
      1 kymus
      2 kynologisch
      2 kynurenin
      5 kynurensyra
      1 kyoga
      1 kyogá
      1 kyphosis
      1 kyrett
      1 kyrka
     25 kyrkan
     14 kyrkans
      1 kyrkböcker
      1 kyrkby
      2 kyrklig
      2 kyrkliga
      2 kyrkoböcker
      1 kyrkobyggnader
      1 kyrkodörren
      1 kyrkogård
      1 kyrkogårdar
      1 kyrkogården
      1 kyrkoledare
      1 kyrkomålning
      3 kyrkor
      1 kyrkorna
      1 kyrkostaten
      2 kyrkotukt
      1 kyrkotukten
      1 kysk
      1 kyska
      7 kyskhet
      1 kyskhetsbälte
      5 kyskhetsbälten
      1 kyskhetsbältet
      1 kyskhetsbuden
      6 kyssar
      1 kyssjuka
     20 l
      8 la
      1 labans
      2 labarraque
      1 labbprover
      1 labckonceptet
      1 laberinto
      1 labetalol
      1 labia
      1 labial
      1 labiala
      1 labil
      1 labilis
      1 labilitet
      1 lablab
      1 lablistan
      1 labor
      1 laboratorieanalyser
      3 laboratoriebruk
      1 laboratoriedirektören
      2 laboratorieförsök
      2 laboratorieinstrument
      2 laboratoriemiljö
      1 laboratorieolyckor
      2 laboratorieprov
      1 laboratorieprover
      6 laboratorier
      1 laboratories
      2 laboratoriestudier
      3 laboratoriet
      2 laboratorietest
      8 laboratorietester
      1 laboratorietesterna
      1 laboratorieundersökning
      1 laboratorieundersökningar
      3 laboratorieutrustning
      1 laboratorieutvärderingar
      1 laboratorieverifierades
      1 laboratoriska
     13 laboratorium
      3 laboratory
      1 labour
      2 labprover
      2 labrador
      1 labretpiercingar
      1 labretpiercingen
      3 laburnum
      1 labyrint
      1 labyrinten
      1 lacadémie
      3 lacan
      3 lacaniansk
      4 lacevaran
      1 lachesis
      2 lack
      1 lacka
      2 läcka
     10 läckage
      2 läckande
      2 lacker
     23 läcker
      3 läckt
      1 lacmoid
      1 lactarius
      1 lactea
      1 lactobaccillus
      1 lactobaciller
      2 lactobacillus
      3 lada
      3 låda
      3 lådan
      1 ladda
      7 laddad
      9 laddade
      2 laddar
      5 laddas
      1 laddat
     13 laddning
      2 laddningar
      1 laddningarna
      4 laddningen
      2 laddningsbara
      1 laddninngsbart
     20 lade
     12 läder
      2 läderaktigt
      4 läderartade
      1 läderband
      1 läderetui
      1 läderhandskar
      2 läderhud
      3 läderhuden
      1 läderkängor
      2 läderpåse
      1 läderstrigel
     16 lades
      1 lådor
      2 ladugårdar
      1 ladugården
      1 lady
      1 läekemedel
      1 laesa
      1 laesio
      1 laetiflorus
      1 laetrile
     44 lag
    177 låg
      4 laga
    114 låga
      1 lagade
      1 lågaktiv
      2 lågan
      1 lagändring
      1 lagändringar
      1 lagändringarna
      2 lagändringen
     24 lagar
      1 lagarna
      2 lagberg
      1 lågblad
      1 lågbr
      1 lagd
      1 lagde
      1 lågdensitetslipoproteiner
      1 lågdos
      1 lågdosantibiotika
      1 lågdosbehandling
      1 lågdosdatortomografi
      2 lågdoserat
      2 lågdosstrålning
     33 läge
      2 lågeffektlaser
      1 lågeffektslaser
     31 lagen
      1 lägen
      1 lågenergilampor
      2 lägenheten
      4 lägenheter
      2 lagens
     36 lager
      4 läger
      1 lagerblad
      1 lagercrantz
      1 lagerhägg
      1 lagerhållning
      1 lagerkörsvatten
      2 lägersmål
      1 lagerträd
      1 lagerträdet
      1 lagerträdets
      1 lägesvarierat
      1 lägesyrsel
      6 läget
      1 lagets
      1 lågfärg
      1 lågfettkost
      1 lågfiberkost
      1 lagföra
      3 lagföreskrifter
      1 lagförslag
      1 lågfrekvent
      4 lågfrekventa
      4 lägg
     49 lägga
     17 läggas
      1 läggdags
     60 lägger
      4 läggning
      1 läggningar
      2 läggningen
      1 låggradig
      1 låggradiga
      1 låggradigt
     47 läggs
      3 låginkomstländer
      1 lågintensiv
      1 lågintensivt
      1 lågkalorikost
      1 lågkalorimetoden
      1 lågkolhydradieter
      1 lågkolhydrat
      7 lågkolhydratdiet
      2 lågkolhydratdieter
      1 lågkolhydratkost
      1 lågkolhydratskost
      1 lagkrav
      1 låglaktosmjölk
      7 laglig
      2 lagliga
      1 lagligen
      7 lagligt
      1 laglöshet
      1 laglöst
      2 laglydigt
      1 lågmolekylära
      1 lågmolekylärt
      1 lagning
      7 lagom
      1 lågpresterande
     10 lagra
      1 lagrad
      1 lagrade
      6 lagrar
     17 lagras
      3 lagrat
      1 lagrats
    145 lägre
      1 lagreglerad
      1 lagregleringar
      3 lagren
     13 lagret
      2 lagring
      1 lagringsförmåga
      1 lagringskärlet
      1 lagringsplats
      2 lagringstid
      2 lagringstiden
      2 lågrisk
      1 lågriskvirus
      1 lagrum
      7 lägst
     12 lägsta
      1 lagstadgad
      1 lagstifta
      1 lagstiftades
      1 lagstiftare
     19 lagstiftning
      1 lagstiftningar
      8 lagstiftningen
      1 lagstiftningens
     12 lagt
     75 lågt
      1 lågteknologisk
      1 lagtexten
      1 lågtröskelverksamhet
      1 lågtröskelverksamheter
      5 lagts
      1 lågvarvsborr
      1 lågvarvsborren
      1 lågväxande
      1 lågväxt
      1 lain
      5 laing
     19 läka
      1 lakan
     12 läkande
      1 läkandeprocessen
      2 lakanen
      2 läkar
      1 läkarbedömningar
      7 läkarbesök
    240 läkare
      2 läkared
    108 läkaren
      6 läkarens
      3 läkares
      1 läkaresällskapet
      2 läkaresällskapets
      3 läkarexamen
      2 läkarförbund
      1 läkarförbundet
      2 läkarhjälp
      1 läkarintyg
      5 läkarkåren
      1 läkarkontroller
      1 läkarlatin
      5 läkarlegitimation
      1 läkarlicens
     13 läkarna
      2 läkarnas
      1 läkarrapporter
      1 läkarrättegången
      1 läkarsällskap
      1 läkarspråket
      1 läkarsprit
      1 läkarstation
      1 läkarstudenter
      1 läkartäthet
      1 läkarteamet
     10 läkartidningen
      1 läkartjänst
      5 läkarundersökning
      1 läkarutbildning
      1 läkarutbildningen
      1 läkarutbildningskommitté
      8 läkarvård
      3 läkarvården
      1 läkarverksamhet
      3 läkarvetenskapen
      2 läkarvetenskapens
      3 läkaryrket
      2 lakas
      4 läkas
      3 lake
      1 läkeageratum
      2 läkebok
      1 läkeeurytmi
      4 läkeeurytmin
      1 läkeeurytmins
      1 läkeeurytmiska
      1 läkeguden
      8 läkekonst
      7 läkekonsten
      4 läkekonstens
      1 läkekunige
      1 läkekunnige
      1 läkemdel
    484 läkemedel
      3 läkemedels
      1 läkemedelsanvändning
      1 läkemedelsavdelning
      2 läkemedelsbehandlad
     17 läkemedelsbehandling
      3 läkemedelsbehandlingar
      2 läkemedelsbehandlingen
      1 läkemedelsberedningar
      1 läkemedelsberoende
      3 läkemedelsbiverkning
      4 läkemedelsbiverkningar
      1 läkemedelsboken
      1 läkemedelsbolag
      1 läkemedelsbolaget
      1 läkemedelsbutiker
      1 läkemedelsexanthem
      2 läkemedelsexpert
      1 läkemedelsfakta
     11 läkemedelsföretag
      1 läkemedelsföretagen
      7 läkemedelsföretaget
      1 läkemedelsförmånen
      1 läkemedelsförmånsverket
      1 läkemedelsförsäkringen
      1 läkemedelsgenomgångar
      1 läkemedelsgivning
      2 läkemedelsgrupp
      1 läkemedelsgrupper
      1 läkemedelsguiden
      1 läkemedelshistorien
      6 läkemedelsindustrin
      1 läkemedelsintag
      2 läkemedelskandidater
      2 läkemedelskemi
      2 läkemedelsklass
      1 läkemedelsklassen
      1 läkemedelsklasser
      1 läkemedelsklassning
      1 läkemedelskombinationer
      1 läkemedelskontroll
      1 läkemedelskostnader
      1 läkemedelsmetaboliter
      1 läkemedelsmissbrukare
      2 läkemedelsmyndigheten
      1 läkemedelsnamnet
      1 läkemedelsområdet
      3 läkemedelsöverkänslighet
      1 läkemedelsprodukt
      1 läkemedelsprodukter
      1 läkemedelsprövning
      2 läkemedelsreaktioner
      1 läkemedelsrelaterade
      2 läkemedelsresistenta
      1 läkemedelsstudier
      4 läkemedelssubstans
      1 läkemedelssubstansen
      3 läkemedelssubstanser
      1 läkemedelssyntes
      2 läkemedelsterapi
      1 läkemedelstillverkning
      1 läkemedelstyperna
      1 läkemedelsupplysning
      1 läkemedelsurval
      1 läkemedelsutlösta
      1 läkemedelsvärderingar
     31 läkemedelsverket
      6 läkemedelsverkets
      1 läkemedelverket
     32 läkemedlen
      1 läkemedlens
     55 läkemedlet
      5 läkemedlets
      1 [läke]ört
      1 läkeprocess
      3 läkeprocessen
      1 läkeprocesser
     22 läker
      1 läkesprocessens
      1 läketiden
      1 läkeväxt
      2 läkeväxten
      1 läkeväxter
      1 lakning
     15 läkning
     12 läkningen
      1 läkningsförmåga
      1 läkningsprocess
      1 läkningsprocessen
      2 läkningsprocesser
      1 lakrits
      1 läks
     10 läkt
      3 läkta
      1 laktamantibiotika
      1 laktamringen
      9 laktas
      1 laktasbrist
      2 laktasenzym
      2 laktaset
      1 laktasgenens
      1 laktasnivåer
      1 laktastabletter
      9 laktat
      3 laktatacidos
      4 laktatdehydrogenas
      1 laktatet
      1 laktationen
      1 laktationens
      1 laktationspsykos
      1 laktatnivåerna
      1 laktatstrukturen
      1 lakterande
      1 läktiden
      1 laktobaciller
      1 lakton
      1 laktoovovegetarianer
     21 laktos
      1 laktosbaciller
      5 laktosen
      2 laktosfri
      1 laktosfria
      1 laktosinnehåll
     25 laktosintolerans
      2 laktosintolerant
      6 laktosintoleranta
      1 laktosnivån
      1 laktostoleranta
      1 laktovegetarianer
      1 laktulos
      1 lalein
      2 lalia
      1 lalía
      1 lambanein
      2 lambda
      1 lamberteatons
      1 lamblia
      1 lameller
      1 lamellerat
      3 lamellerna
      1 lamfetamin
      1 lamictal
      9 lamin
      5 lamina
      1 laminat
      1 laminer
      1 lamingenen
      1 laminin
      1 lämlar
      4 lamm
     30 lämna
      8 lämnade
      4 lämnades
      4 lämnande
     33 lämnar
     22 lämnas
      6 lämnat
      4 lämnats
      2 lämningar
      1 lämningarna
     10 lampa
      2 lämpad
      4 lämpade
      3 lampan
      1 lampans
     16 lämpar
      1 lampglaset
     40 lämplig
     24 lämpliga
      2 lämpligare
      2 lämpligast
      2 lämpligaste
      3 lämplighetstest
     25 lämpligt
      1 lampor
      1 lamprocapnos
      1 lån
     32 län
      6 låna
      1 lånade
      2 lånades
      2 lånar
      1 lånat
      1 lånats
      1 lanceolata
     10 lancet
      1 lanc�me
     34 land
      6 landar
      1 landat
      1 landehag
    367 länder
      1 länderm
     23 länderna
      1 ländernas
      9 länders
     52 landet
      9 landets
      1 landis
      2 ländkota
      1 ländkotan
      1 ländkotorna
      1 landkrokodil
      1 landkrokodilen
      2 landlevande
      1 landmärke
      1 landormar
      7 ländryggen
      1 ländryggsbesvär
      1 ländryggsmärta
      2 ländryggssmärta
      3 lands
      1 landsända
      1 landsbygd
     10 landsbygden
      2 landsbygdens
      1 landsbygdskommuner
      2 landsbygdsområden
      1 landsflyktiga
      1 landskapsblomma
      1 landskapslagarna
      1 landskapssvamp
      1 landsknekt
      1 landsköldpaddor
      1 landskontor
      1 landsnäcka
      2 landsortspolis
      1 landsortssjukhusen
      4 landsteiner
     23 landsting
     10 landstingen
      3 landstingens
      1 landstinges
      4 landstinget
      1 landstingets
      1 landstingsfullmäktige
      1 landstingskommunal
      1 landväxter
      1 landvinningar
      1 landyta
      1 lane
      1 lånemöjligheter
      1 lånemöjligheterna
      1 länenslandstingens
      1 lånereglerna
      2 länet
      1 lanfranc
      1 lang
    181 lång
    114 långa
      1 långärmad
      1 långbågar
      2 långbåge
      1 långbyxor
     44 längd
      1 längdavstånd
     23 längden
      2 längder
      2 långdistanslöpare
      2 långdragen
      1 långdragenhet
      2 långdraget
      2 långdragna
      1 längdriktning
      1 längdskidåkning
      2 längdtillväxt
    148 länge
      1 langerhanscell
      6 langerhanska
      1 långfibrig
      1 långfilmen
      1 långfingret
      1 långivare
      1 långkedjig
      1 långkörningar
      1 långlivad
      4 långlivade
      1 långlivat
      1 langogne
      1 långpromenader
    292 längre
      1 långresa
      1 långresor
      3 langs
     55 längs
     26 långsam
      2 långsamhet
     12 långsamma
     22 långsammare
     57 långsamt
      1 långsamväxande
      1 långsegling
      1 långsele
      3 längsgående
      7 långsiktig
     12 långsiktiga
     10 långsiktigt
      2 långsiktligt
      2 långskaftade
      1 långskalle
      1 långsmal
      1 långsmala
     22 längst
      8 längsta
      1 långsträckta
    125 långt
      3 längtan
      1 långtgående
      1 långtida
      1 långtidsanvändning
      1 långtidsbehandling
      1 långtidsbehandlingar
      1 långtidseffekt
      1 långtidseffekter
      2 långtidsminne
      1 långtidsresultat
      1 långtidssmittade
      3 långtidsstudier
      1 långtidsuppföljning
      1 långtidsuppföljningar
      1 långtidsuppföljningsstudier
      1 långtidsutkomst
      1 långtidsutövare
      1 långtidsverkan
      3 långtidsverkande
      1 långväga
      1 långvård
     84 långvarig
     31 långvariga
      1 långvarigare
     27 långvarigt
      4 långverkande
      1 langworthy
      7 länk
      2 lanka
      1 länkad
      2 länkade
      1 länkadt
     27 länkar
      1 länkas
      1 länkat
      3 länken
      1 länkning
      1 la�nnec
      3 lånord
      3 lånordet
      1 lans
      4 läns
      1 länsdelssjukhus
      2 lansera
      1 lanserad
     11 lanserade
     18 lanserades
      2 lanseras
      1 lanserat
      7 lanserats
      1 lansering
      3 lanseringen
      2 lansett
      1 lansettapparat
      1 lansetter
      2 lansettfiskar
      1 lansettfönster
      4 lansettlika
      2 länslasarett
      1 lanslika
      1 länsrätten
      1 länsstyrelse
      1 länsstyrelsernas
      1 lanszwertii
      1 lantbor
      1 lantbrukare
      1 lantbrukarna
      1 lantbruket
      1 lantbruksdjur
      1 lantbruksspruta
      2 lantbruksuniversitet
      1 lantern
      1 lantmannen
      1 lantmäteri
      1 lantus
      1 lanzoprazol
      1 lapa
      1 laparoskop
      1 laparoskopet
      1 laparoskopi
      2 laparoskopisk
      1 laparotomi
      1 laparotomier
      1 lapis
      1 lapisdroppar
      1 lapp
      4 läpp
     18 läppar
     17 läpparna
      2 läpparnas
      5 läppbalsam
      1 läppbalsamläppcerat
      1 läppcerat
      1 läppcyanos
      5 läppen
      3 läppförstoring
      1 läppiercingarna
      1 läppiercingen
      2 lappland
      1 läpplattor
      1 läpppiercing
      1 läpppiercingar
      1 läpppiercingen
      1 läppsmycket
      8 läppstift
      3 läpptallrikar
      1 lapraskopi
      1 lapraskopiska
      1 lapraskopiskt
      6 lår
     18 lär
      1 lara
     47 lära
     53 läran
      8 lärande
      3 lärandet
      1 lärans
     15 lärare
      1 lärarpåverkan
      1 läras
      2 lårben
      2 lårbenet
      1 lårbenets
      1 lärda
      8 lärde
      1 lärdes
      1 lärdomarna
      4 låren
      1 lårens
      3 låret
      1 lårets
      1 lårficka
      1 lariam
      4 lärjungar
      2 lärjunge
      1 lärjungeförhållande
      2 lärling
      1 lärlingens
      1 lärlingstiden
      5 larm
      1 larmarmband
      1 larmas
      1 larmen
      3 larmet
      1 larmläkemedel
      1 larmnummer
      1 larmrapporter
      2 larmsignaler
      1 larmstation
      2 larmtjänst
      4 läroböcker
      1 läroplan
      1 läror
      1 lärosäten
      1 lärosätena
      1 lärosätets
      1 lärosatser
      1 larry
      8 lars
      1 lärs
      1 larsen
      1 larserik
      1 larsgöran
      1 larsgunnar
      2 larsson
     11 lärt
      7 larv
      1 larvartad
      1 larvbenämningarna
      8 larven
     34 larver
     33 larverna
      1 larvformer
      1 larvstadier
      2 larvstadiet
      5 laryngektomi
      2 laryngit
      1 laryngofarynx
      1 laryngopharynx
      3 laryngoskop
      2 laryngoskopet
      2 laryngospasm
      4 larynx
      3 las
      1 lås
     24 läs
      4 låsa
     38 läsa
      2 läsande
      1 läsandet
      1 låsanordning
      1 läsare
      2 läsaren
      1 läsarens
      1 läsåret
     14 lasarett
      3 lasaretten
      1 lasarettsläkare
      1 lasarettsstadgans
      1 läsas
      1 låsbar
      1 lascaux
     16 laser
      3 låser
      6 läser
      4 laserbehandling
      1 laserdopplerteknik
      1 laserfibrer
      1 laserkateter
      1 laserkirurgi
      1 laserkirurgin
      1 laserklass
      2 laserljus
      1 laserljuset
      3 lasern
      2 laserstråle
      4 laserterapi
      3 läses
      1 läsflyt
      2 läsförmåga
      1 läsförmågan
      1 läsförståelsen
      1 läsfunktionen
      1 läsglasögon
      1 läshandikapp
      1 läshinder
      1 läsinlärningen
      1 lasix
      2 läsk
      2 läskedrycker
      4 lasker
      4 laskerpriset
      1 laskerstiftelsen
      1 läskpappersbitar
      1 läskpappret
      1 läskunniga
     15 läsning
      1 läsningar
      7 läsningen
      1 läsningsfel
      1 låsningsfria
      1 läspning
      1 läsproblem
      2 lasrar
      1 läsrelaterade
      1 lassa
     12 lassafeber
      2 lassavirus
      1 lasset
      2 lassonde
      1 lässvårighet
      7 läst
      1 låsta
      1 lästa
      1 lastade
      1 lastbärande
      1 lastbilar
      1 lastbilschaufförer
      3 läste
      2 lasten
      1 lästes
      1 lästilläggets
      1 läsuttal
      1 läsverktyg
     25 lat
      6 låt
     10 lät
      1 lata
     47 låta
      1 latah
      2 låtar
      1 låtarna
      1 latensintervallet
      1 latenstiden
      1 latensvariationer
     31 latent
      4 latenta
     41 låter
      2 lateral
      5 laterala
      1 lateralis
      1 lateralt
      9 latex
      1 latexagglutinationstest
      1 latexallegiker
      1 latexallergiker
      2 latexen
      2 latexkatetrar
      1 latexkondom
      1 latexöverkänslig
      2 lathyrism
    134 lathyrus
     88 latin
      3 latinamerika
      1 latinamerikaner
      2 latinamerikansk
      2 latinet
     39 latinets
      2 latinisering
      1 latinsk
     24 latinska
      4 latinskt
      5 låtit
      1 latituderna
      1 låtna
      1 latrin
      2 låtsas
      1 lått
    147 lätt
     24 lätta
      1 lättade
      1 lättantändlig
      1 lättantändliga
      1 lättantändlighet
      2 lättantändligt
      2 lättanvänt
      2 lättar
      2 lättarbetad
    104 lättare
      6 lättast
      4 lättaste
      1 lättat
      1 lättåtkomliga
      1 lättbearbetad
      1 lättbearbetade
      1 lättbehandlade
      1 lättdistraherad
      1 lättfattlig
      2 lättflyktig
      1 lättflyktiga
      1 lättflyktighet
      2 lättflytande
      1 lättförklarlig
      1 lättförståeliga
      2 lätthanterliga
      1 lätthanterligt
      1 lätthet
      1 lättigenkännliga
      1 lättillgänglig
      1 lättillverkat
      1 lättja
      1 lättjusterade
      1 lättkammat
      1 lättkritiserad
      3 lättlöslig
      3 lättlösliga
      4 lättlösligt
      1 lättmetall
      2 lättmetaller
      3 lättnad
      3 lättnadskänsla
      2 lättodlad
      1 lättoxiderade
      2 lättretlighet
      1 lättrinnande
      2 lättskött
      1 lättsmältt
      1 lättstyrd
      1 lättvårdsgruppen
      1 lättviktiga
      1 lättvindig
      1 latum
      2 laudanum
      2 laura
      1 laurent
      1 laurocerasi
      1 laurocerasin
      1 laurocerasus
      2 lav
      1 lavabo
      1 lavar
      1 lavarna
      1 lavely
     22 lavemang
      3 lavemanget
      1 lavemangstillsats
      1 laven
      1 lavendel
      1 lavoisier
      1 law
      1 lawford
      3 lawrence
      2 lax
      1 läxa
      1 laxantia
      2 laxativ
      1 laxativa
      1 laxer
      2 laxerande
      2 laxering
      5 laxermedel
      1 laxfärgade
      1 laxiflorus
      1 läxor
      1 laxrosa
      1 layardii
      1 layout
      1 lazareth
      1 lazzaretto
      1 lbp
      1 lcdskärm
      4 lchf
      1 lchfdieter
      1 lchfförespråkare
      1 lchfmetoden
      1 lcmv
     10 ld
      1 ldalocal
      2 ldd
      1 lddosen
      4 ldh
      3 ldl
      7 ldlkolesterol
      1 ldopa
      1 ldvärde
      5 le
      1 leaf
      1 league
      1 learn
      1 least
      1 lebensborn
      2 lebensbornkliniker
      1 lebensbornprogrammet
      2 leber
      1 leberecht
      1 lecitin
      1 leclaire
      1 lectin
      5 lectularius
     56 led
    350 leda
      1 ledade
      1 ledamoten
      2 ledamöter
     23 ledande
     10 ledare
      5 ledaren
      1 ledarforum
      6 ledarhund
     10 ledarhundar
      7 ledarhunden
      1 ledarhundens
      1 ledarhundsdagen
      1 ledarhundsförare
      2 ledarhundsföraren
      1 ledarskap
      1 ledas
      2 ledband
      1 ledbandet
      6 ledbesvär
      1 ledbesvären
      1 ledbrosk
      4 ledbrosket
      4 ledd
      1 ledda
     56 ledde
      2 leddes
      1 leddestruktion
      1 leddjur
      1 ledebouri
     13 leden
      1 ledens
    498 leder
     13 lederna
      1 leders
      4 ledet
      1 ledford
      1 ledförslitning
      1 ledfunktionen
      1 ledgångs
      7 ledgångsreumatism
      1 ledhinnorna
      2 ledi
      2 ledig
      1 ledighet
      2 ledigt
      1 ledinfektioner
     10 ledinflammation
      2 ledinflammationer
      1 ledkapsel
      2 ledkapslar
      1 ledkula
      9 ledning
      3 ledningar
      1 ledningarna
      2 ledningen
      1 ledningsansvariga
      1 ledningsbana
      2 ledningsbanan
      1 ledningsbanorna
      1 ledningsbunden
      1 ledningsfibrerna
      2 ledningsförmåga
      2 ledningshastighet
      1 ledningsnät
      1 ledningsnäten
      1 ledningssträckor
      2 ledningssystem
      1 ledpanna
      1 ledprotes
      2 ledproteser
      1 ledpunktion
     16 leds
      2 ledsamhet
      1 ledsamma
      5 ledsen
      1 ledsjukdom
      3 ledsjukdomar
      1 ledsmärtor
      1 ledsvullnad
      7 ledtrådar
      1 leduc
     11 ledvärk
      2 ledvätska
      1 ledvätskor
      2 ledvätskorna
      1 ledverk
      1 ledytan
      1 ledytorna
      4 lee
      1 leem
      3 leende
      1 leeuwenhock
      3 leeuwenhoek
      2 legal
      6 legala
      1 legalförskrivning
      1 legalisera
      1 legaliserat
      1 legalisering
      1 legalitet
      1 legalt
      9 legat
      2 legend
      1 legendarisk
      1 legenden
      1 legender
      1 legerat
      6 legering
      2 legeringar
      1 legion
      6 legionärssjuka
      1 legionärssjukan
     14 legionella
      1 legionellaarter
      2 legionellabakterien
      2 legionellabakterier
      1 legionellabakterierna
      1 legionellaceae
      1 legionellaproblem
      1 legionellautbrott
      2 legionellautbrotten
      1 legislativt
      1 legitim
     23 legitimation
      1 legitimationen
      1 legitimationer
      3 legitimationsgrundande
      1 legitimationsyrke
      2 legitimera
     15 legitimerad
     20 legitimerade
      1 legitimerande
      1 legitimerar
      2 legitimerat
      1 legitimitet
      2 legitimt
      1 legosoldat
      2 legosoldater
     10 lehmann
      2 lehmanns
      1 lehrbuch
      2 leibniz
      1 leiden
      3 leif
      1 leijonborg
      1 leiomyom
      7 leiomyosarkom
      1 leipzig
      1 leishmaniasis
      1 lejon
      1 lejonansikte
      1 lejonparten
      1 lejour
      8 lek
      1 leka
      1 lekande
      2 lekar
      2 lekartävlingar
      1 leken
      3 leker
      1 lekhjälm
      2 lekman
      7 lekmän
      2 lekplatser
      1 leksaker
      2 leksell
      1 lekte
      2 lektiner
      1 lem
      1 lemförlängningskirurgi
      7 lemmar
      1 lemmarna
      2 lemmen
      1 lemmissbildningar
      1 lena
      1 lenande
      1 lengberg
      1 lennart
      2 lennon
      1 lennonplastic
      2 lenny
      1 lentiformis
      1 lentinus
      1 lentis
      1 lentivirus
      2 lenvironnement
      1 leo
      6 leonard
      4 leonardo
      4 leone
     19 lepra
      1 leprabakterien
      4 leprae
      1 leprakolonier
      1 leprapatienter
      2 leprasjuka
      2 lepromatösa
      1 lepromatosis
      1 leprosarium
      1 lepsis
      4 leptin
      2 leptosphaeria
      5 leptospiros
      2 ler
      3 lera
      1 lerfigur
      1 lergigan
      1 lergods
      1 lerjord
      1 lermark
      2 leror
      1 lerplattor
      1 lerskreppe
      1 lertavlor
      1 les
      3 lesion
      2 lesionen
      7 lesioner
      2 lesionerna
      8 leta
      3 letade
      1 letades
      3 letal
      2 letala
      3 letalitet
      2 letaliteten
      1 letandet
     12 letar
      2 letargi
      2 letat
      2 lethal
      1 letrozol
     47 lett
      1 letter
      1 letterbyletter
      1 letters
      1 lettiskans
      1 lettland
      1 leucanthus
      9 leucism
      1 leucistisk
      2 leucistiska
      1 leucistiskt
      1 leuckarts
      1 leucokori
     28 leukemi
      4 leukemier
      2 leukemipatienter
      1 leukemoid
      1 leukocyte
     10 leukocyter
      1 leukocyterna
      1 leukocytesteras
      2 leukocytos
      1 leukodermi
      3 leukopeni
      1 leukotil
      1 leukotrienantagonist
      1 leukotrienantagonister
      1 leukotriener
     56 leva
    110 levande
      1 levandefödande
      1 levandefödare
      1 levandefoder
      1 levas
      1 levat
      1 levaxin
     24 levde
      4 level
      1 levels
    154 lever
      1 leveråkommor
      2 leverans
      1 leveransavtal
      3 leveransen
      1 leverantör
      3 leverantörer
      1 leverantörsberoende
      1 leverantörsföreningen
      2 leverbiopsi
      7 levercancer
      3 leverceller
      4 levercellerna
      5 levercirros
      1 leverelastografi
      1 leverencefalopati
      1 leverencefalopatin
      1 leverenzym
      2 leverenzymer
      7 leverera
      1 levererade
      7 levererar
     10 levereras
      1 levererat
      2 levererats
      1 leverereras
      1 leverfläck
      1 leverfläckar
      1 leverfliken
      1 leverflundran
      1 leverflundrans
      1 leverflundror
      1 leverförstoring
      5 leverfunktion
      1 leverfunktionen
      1 leverfunktionsprov
      1 leverfunktionstester
      1 levergång
      2 levergången
      1 leverincision
      1 leverinflammaion
     10 leverinflammation
      1 leverinsufficiens
      1 leverkanten
      3 leverkoma
    134 levern
      3 leverne
      1 levernekros
      8 leverns
      1 leverparasiter
      3 leverpåverkan
      1 leverproblem
      1 leverprover
      1 leversegment
      8 leversjukdom
      6 leversjukdomar
      7 leverskada
     11 leverskador
      1 leverskadorna
      1 leverstärkelse
      2 leverstatus
      1 leverstigmata
      5 leversvikt
      1 levertestvärden
      3 levertransplantation
      1 levertransplantationen
      4 levervärden
      2 levervärdena
      1 levervävnaden
      1 levetiracetam
      1 levin
      3 levines
      1 levitra
      4 levnad
      2 levnaden
      1 levnadsålder
      7 levnadsår
      3 levnadsåren
      5 levnadsåret
      1 levnadsbetingelser
      2 levnadscykel
      1 levnadsdagar
      1 levnadsdygnen
      1 levnadsförhållandena
      1 levnadsmånaderna
      2 levnadsmiljö
      1 levnadsmiljön
      5 levnadsmönster
      1 levnadsnivå
      1 levnadsregler
      1 levnadsreglerna
      7 levnadssätt
      1 levnadsstadier
      2 levnadsstandard
      2 levnadstid
      2 levnadsvanor
      1 levnadsveckor
      3 levnadsvillkor
      4 levoamfetamin
      1 levoamfetaminet
      1 levra
      3 levrar
      1 levras
      1 levrets
      2 levs
     10 levt
      1 lewins
      2 lewis
      1 lewy
      3 lewykroppar
      2 lewykroppatienter
      3 lewykroppsdemens
      2 lex
      1 lexikon
      1 lexis
      4 leydigceller
      3 lformen
      1 lga
      1 lgd
      1 lge
      2 lgg
      2 lglukos
      1 lglutamin
      1 lgm
      8 lh
      1 lhasa
      1 lhrh
      1 lhyoscyamin
      2 liaisonkontor
      1 lian
      1 libani
      1 liber
      2 liberal
      1 liberalisering
      1 liberaliseringens
      3 liberia
      1 libertarianism
      1 liberties
      9 libido
      1 [libido]
      2 libidon
      6 libidot
      2 libidots
      1 libra
      2 libresse
      2 lice
      5 licens
      1 licensbelagda
      1 licensierade
      1 licensinnehavaren
      1 licenstvånget
     26 lida
     31 lidande
      4 lidanden
      7 lidandet
      1 lidandets
      1 lidcombe
    126 lider
      2 lidingö
      5 lidit
      2 lidokain
      1 liebig
      1 liechtenstein
      1 lien
     10 life
      1 lifestyle
      1 lifta
      2 liftar
      1 liftarens
      1 liftning
      1 lifvet
      1 liga
      5 ligament
      1 ligand
      1 ligandbindning
      1 liganden
      1 ligander
      3 li�ge
      2 ligering
     56 ligga
     21 liggande
    212 ligger
      2 liggsår
      1 lightheadedness
      1 lighting
      1 ligistsubkulturer
      1 lignieresii
      1 lignin
      1 ligninbevarande
      1 ligninet
      8 lik
    197 lika
      1 likabetydande
      7 likadan
      4 likadana
      2 likadant
      7 likaledes
      1 likande
      1 likaregeln
      6 likartad
     10 likartade
      2 likartat
     35 likaså
      2 likaväl
      1 likbesiktning
      1 likblå
      3 like
      3 liket
      1 likgift
      4 likgiltighet
     34 likhet
      4 likheten
     16 likheter
      1 likheterna
      1 likkall
      1 likkörarna
     20 likna
      7 liknade
    217 liknande
     87 liknar
     16 liknas
      1 liknelsen
      1 liko
      1 liköppningar
      1 likörtillverkning
      1 likrikta
      1 likriktning
      1 liksidig
      1 liksidigt
    147 liksom
      1 likspänning
      1 likspänningskomponenter
      1 likställa
      1 likställas
      2 likställda
      2 likställdes
      1 likställigt
      1 likställs
      3 likström
     25 likt
      1 liktornar
      1 liktydig
      2 liktydigt
      9 likväl
      3 likvärdig
      4 likvärdiga
      3 likvärdigt
      1 likvärt
      2 likvor
      1 likvorprover
      4 lila
      1 lilaaktiga
      1 lilablå
      1 liliaceae
      1 liliales
      2 lilium
      1 lilja
      3 liljekonvalj
      2 liljekonvaljen
      2 liljekonvaljens
      1 liljekonvaljer
      1 liljekonvaljerna
      1 liljesläktet
      3 liljeväxter
      3 liljeväxterna
     18 lilla
      1 lille
      1 lillfinger
      1 lillfingret
      1 lillhjärna
      6 lillhjärnan
      3 lilltå
      1 lilltåa
      2 lilltån
      1 lim
     11 limbiska
      2 lime
      1 limejuice
      1 limey
      1 limfilmen
      2 limited
      1 limma
      1 limmade
      1 limmet
      2 limning
      1 limnologi
      5 limonen
      1 limulus
      8 lin
      1 linac
      1 linalool
      1 linamarin
      1 linan
      6 lind
      3 linda
      1 lindad
      1 lindar
      1 linde
      1 linderefref
      1 lindgrens
      1 lindning
     56 lindra
      1 lindrade
      1 lindrades
      4 lindrande
     14 lindrar
     12 lindras
     18 lindrig
     12 lindriga
     30 lindrigare
      1 lindrigast
      1 lindrigaste
      6 lindrigt
     10 lindring
      1 lindsay
      1 lindström
      6 linea
      2 linear
      1 linearifolius
      2 linezolid
      3 linfrö
      1 linfrön
      2 linfröolja
      1 ling
      1 lingam
      1 lingua
      8 linguae
      1 lingual
      1 linguala
      2 lingvistik
      1 lingvistisk
      1 linifolius
      2 liniment
      2 linjaler
      5 linjär
      1 linjära
      1 linjäraccelerator
      1 linjäracceleratorer
      3 linjäracceleratorn
      6 linjärt
     12 linje
      6 linjen
     11 linjer
      3 linjerna
      1 linjespecifika
     11 linköping
      4 linköpings
      1 linkosamider
      8 linne
     10 linné
      1 linnen
      1 linnepressen
      1 linnés
      2 linnet
      1 linnetyg
      2 linnéuniversitetet
      1 linnevaror
      1 linnevarorna
      1 linoleic
      1 linolensyra
      1 linoleummattor
      1 linolsyra
      2 linor
     12 lins
      1 linsanvändning
      1 linsbärare
      1 linsbevarande
     14 linsen
      7 linsens
     21 linser
     11 linserna
      1 linskapseln
      1 linskolobomoch
      3 linsluxation
      1 linsmarknaden
      1 linstyp
      1 linstyper
      1 linsvätska
      1 lintyg
      1 lionizes
      1 lipanthyl
      4 lipas
      2 lipaser
      2 lipid
      1 lipiddel
      1 lipiddelen
      4 lipider
      2 lipidhölje
      1 lipidhöljen
      1 lipidlager
      1 lipidstruktur
      3 lipitor
      1 lipo
      1 lipodermatoscleros
      1 lipodystrofi
      4 lipolys
      5 lipom
      2 lipomet
      1 lipomyelomeningocele
      1 lipooligosackarider
      1 lipopolysackarid
      3 lipopolysackarider
      2 lipoprotein
      2 lipoproteiner
      1 lipoproteinlipas
      1 lipoptena
      2 liposarcom
      1 liposarkom
      4 liposom
      1 liposomen
      4 liposomer
      1 liposomerna
      1 liposuction
      1 lipoteichoic
      1 lipoteikonsyra
      1 lipskys
      1 liquide
      1 liquor
      1 lirka
      1 lirkas
      2 lisdexamfetamindimesylat
      1 lisdexamfetamindimesylatet
      1 lisn
      1 lissajouskurvor
      2 list
     20 lista
      2 listad
      5 listade
      1 listades
      4 listan
      3 listar
     10 listas
      1 listats
      3 listen
      1 listeria
      1 listeriaförgiftning
      1 listerios
      1 listers
      1 listor
      1 lita
      1 litauen
      1 litauenfödda
    115 lite
    150 liten
      1 litenhet
     23 liter
      1 literacy
      1 litermin
      1 literminut
      1 liters
      1 litersekund
     60 litet
      1 litharge
      1 lithium
      1 lithopedion
      1 lithopedioner
      1 lithopone
      2 lithos
      4 litium
      1 litterär
      3 litterära
      1 litterärt
     34 litteratur
     28 litteraturen
      1 litteraturens
      1 litteraturgenomgång
      1 litteraturhistoriens
      6 litteraturöversikt
      1 litteraturöversikter
      1 litteraturterapi
      1 little
      1 littoralis
      1 litvinenko
    198 liv
      1 livbåtar
      1 livbåtsfot
      1 livedo
      1 livegna
      1 liver
      1 liverpool
      1 livestocks
    132 livet
      1 livet[]
      1 livetbr
     20 livets
      1 livförsäkring
      1 livförsäkringen
      1 livgarde
      2 livgivande
      1 livhanken
      1 livingstone
      1 livkärnfrisk
      1 livläkare
      1 livläkaren
      2 livlig
      1 livligt
      1 livmedicus
     20 livmoder
      1 livmodercancer
      2 livmoderframfall
      1 livmoderhålan
      2 livmoderhals
     14 livmoderhalscancer
     23 livmoderhalsen
      1 livmoderhalsgångens
      3 livmoderhalskanalen
      1 livmoderhalssekretet
      1 livmoderinflammation
      2 livmoderinnehållet
      4 livmodermunnen
     80 livmodern
      8 livmoderns
      1 livmoderruptur
      2 livmoderscancer
      3 livmoderslemhinna
     11 livmoderslemhinnan
      1 livmoderstappen
      1 livmoderstorlek
      1 livmoderstrakten
      4 livmodertappen
      1 livmodertrakten
      3 livmoderväggen
      1 livmodervävnaden
      9 livnär
      1 livnärt
      1 livomständigheter
      2 livräddande
      2 livräddning
      1 livre
      1 livrem
      1 livs
      1 livsår
      1 livsåskådningar
      2 livsblad
      1 livschanser
     20 livscykel
      3 livscykeln
      1 livsdrift
      3 livsdugliga
      1 livsdugligt
      1 livsdyrkan
      4 livsenergi
      1 livsenergier
      1 livserfarenheter
      1 livsfara
      1 livsfaran
      2 livsfarlig
      2 livsfarliga
      2 livsfarligt
      1 livsförhållanden
      5 livsföring
      2 livsföringen
      1 livsformer
      1 livsfrukt
      1 livshållning
      1 livshändelse
      3 livshändelser
      1 livshjul
     50 livshotande
      1 livshunger
      2 livsinstinkterna
      9 livskraft
      3 livskraften
      1 livskrafter
      1 livskraftig
      1 livskris
      1 livskriser
      1 livskvalité
      1 livskvalitén
      8 livskvalitet
      3 livskvaliteten
     25 livslång
      3 livslånga
     13 livslängd
     11 livslängden
      1 livslängdsförväntan
      5 livslångt
      1 livsleda
     91 livsmedel
      1 livsmedels
      1 livsmedelsaffären
      4 livsmedelsaffärer
      1 livsmedelsbehov
      2 livsmedelsbistånd
      1 livsmedelsbranchens
      2 livsmedelsburen
      2 livsmedelsburna
      2 livsmedelsbutiker
      1 livsmedelsbutikerna
      1 livsmedelsfabriker
      1 livsmedelsfärgämne
      1 livsmedelsfärgämnen
      1 livsmedelshantering
      1 livsmedelshjälp
      1 livsmedelshygien
      1 livsmedelsindustrier
      2 livsmedelsindustrin
      1 livsmedelskedjan
      1 livsmedelsmikrobiologi
      1 livsmedelsorgan
      3 livsmedelsproducerande
      3 livsmedelsprodukter
      1 livsmedelsproduktionen
      1 livsmedelsprogram
      7 livsmedelstillsats
      1 livsmedelstillsatsen
      1 livsmedelstillsatser
     11 livsmedelsverket
      1 livsmedelsvetenskap
      2 livsmedlen
      7 livsmedlet
      2 livsmedlets
      2 livsmiljö
      1 livsmiljöer
      2 livsmönster
      1 livsnivå
      2 livsnödvändig
      4 livsnödvändiga
      1 livsnödvändighet
      1 livsnödvändigt
      5 livsomständigheter
      1 livsomstörtande
      2 livsprocesser
      1 livsprojekt
      5 livssituation
      3 livssituationen
     23 livsstil
      3 livsstilen
      1 livsstilens
      1 livsstils
      1 livsstilsbetingade
      3 livsstilsfaktor
      4 livsstilsfaktorer
      1 livsstilsförändring
      4 livsstilsförändringar
      1 livsstilsorsaker
      1 livsstilsrelaterat
      1 livssynvinkel
      4 livstecken
     13 livstid
      1 livstiden
      2 livstider
      1 livstids
      3 livstidsprevalens
      6 livstidsprevalensen
      1 livstidsrisk
      1 livstråden
      1 livstycke
      2 livstycket
      1 livsval
      1 livsvatten
      1 livsvetenskaperna
      2 livsviktig
      1 livsviktiga
      3 livsviktigt
      1 livsvillkor
      1 livsvillkoren
      2 livvakt
      2 livvakter
      1 livvaktsorganisationer
      1 livvaktsstyrka
      1 livvaktsstyrkor
      1 liza
      1 lizard
    155 ljud
      1 ljudabsorbenter
      1 ljudabsorberande
      1 ljudanläggning
      1 ljudbaserade
      1 ljudbild
      1 ljudbildande
      1 ljudbilden
      1 ljudbildning
      1 ljudböckerna
      1 ljuddämpande
      1 ljuddämpare
     11 ljuden
      1 ljudenmålet
      1 ljudenoljuden
     44 ljudet
      5 ljudets
      1 ljudeurytmi
      1 ljudeurytmin
      1 ljudexponering
      1 ljudfil
      1 ljudfiler
      1 ljudfilerna
      1 ljudfilmen
      1 ljudfobi
      1 ljudförnimmelser
      1 ljudfrekvens
      1 ljudfrekvenser
      1 ljudimpulserna
      2 ljudirritation
      1 ljudisolerande
      6 ljudkälla
      5 ljudkällan
      3 ljudkänslighet
      1 ljudkänsligheten
      1 ljudkonstnärer
      1 ljudkvalitén
      1 ljudlig
      1 ljudliga
      1 ljudljuskänslig
      1 ljudmätare
      1 ljudmiljö
      1 ljudmiljöer
      1 ljudmystik
      1 ljudnära
      9 ljudnivå
      4 ljudnivåer
      8 ljudnivån
      1 ljudnivåvakt
      1 ljudomfång
      1 ljudorienterad
      1 ljudöverkänslig
      3 ljudöverkänsliga
     14 ljudöverkänslighet
      2 ljudöverkänsligheten
      1 ljudproblem
      1 ljudprocessor
      1 ljudproduktionen
      1 ljudsegment
      1 ljudslang
      1 ljudstimulatorer
      3 ljudstimuli
      1 ljudstruktur
      1 ljudstyrka
      2 ljudstyrkan
      1 ljudsystem
      2 ljudterapi
      1 ljudtics
      1 ljudtrauman
      2 ljudtryck
      1 ljudtrycknivåer
      3 ljudtrycksnivå
      1 ljuduppfattning
      3 ljudvågor
      1 ljudvågsvibrationer
      1 ljuga
      2 ljugandet
      3 ljuger
      1 ljummen
      5 ljummet
      5 ljumskar
      8 ljumskarna
      3 ljumskbråck
      3 ljumske
      8 ljumsken
      2 ljumsksvamp
      1 ljunggren
      1 ljungväxter
      1 ljungväxters
     65 ljus
      7 ljusa
      5 ljusare
      1 ljusbehandling
      1 ljusbestrålning
      2 ljusbilden
      1 ljusblåfärgad
      1 ljusblixtar
      1 ljusbox
      1 ljusbrun
      1 ljuseffekt
      1 ljusenergi
     32 ljuset
      1 ljusets
      1 ljusfenomen
      3 ljusförhållanden
      1 ljusgrön
      1 ljusgröna
      1 ljusgul
      1 ljusgula
      1 ljushärdig
      1 ljushet
      1 ljuskaféer
      3 ljuskälla
      1 ljuskällor
      2 ljuskänslig
      5 ljuskänsliga
      3 ljuskänslighet
      3 ljuskänsligt
      1 ljuslåga
      1 ljuslila
      1 ljuspulser
      1 ljuspunkt
      1 ljuspunkten
      1 ljuspunkter
      2 ljusreflex
      1 ljusröda
      1 ljusrosa
      2 ljusrött
      5 ljusrum
      1 ljusseende
      1 ljussignal
      3 ljussken
      1 ljusskygghet
      1 ljusstark
      3 ljusstyrka
      1 ljusstyrkan
     15 ljust
     10 ljusterapi
      1 ljusterapin
      2 ljusterapirum
      1 ljustunnel
      1 ljusvågor
      1 ljusvågslängder
      1 lkg
      3 lkr
      1 lkr]
      1 lkryptor
      1 lkryptorna
      1 l�l
      6 lllt
      1 lm
      1 lmna
      2 lmp
      1 lmpotenser
      1 lnt
      1 lntmodell
      1 lntmodellen
      2 lo
      1 loads
      1 lob
      1 lobak
      7 lobär
      1 lobärt
      1 lobbat
      1 lobbygrupper
      1 lobbyorganisationer
      1 lobbyverksamhet
      1 lobelia
      1 loben
      5 lober
      2 loberna
      1 lobotomerade
      1 lobotomerades
      1 lobotomerande
      1 lobotomeringarna
      8 lobotomi
      4 lobulära
      3 lobuli
      1 lobulus
      1 lobus
      1 locis
      4 lock
      3 locka
      1 lockad
      3 lockande
      8 lockar
      2 lockas
      2 locke
      1 locked
      2 lockedintillstånd
      1 locket
      1 lockets
      1 lockigt
      1 locktänger
      2 locus
      1 lod
      2 löd
      1 löda
      2 lödas
      2 lödder
      1 löddrade
      1 loddrar
      2 löddrar
      1 löddret
      1 löder
      1 lödkolv
      1 lödning
      3 lodräta
      1 lodstrykjärnen
      1 lodstrykjärnet
      1 loe
      1 loftbastun
      1 löfte
      1 löften
      1 loftet
      1 löfven
      1 log
      1 logaritmen
      1 logaritmeras
      1 logaritmform
      1 logaritmisk
      1 logaritmiskt
      1 logaritmlagarna
      1 logho
      1 logia
      1 logik
      2 logikanalysator
      2 logikanalysatorn
      1 logiké
      3 logisk
      1 logiska
      1 logiskmatematisk
      4 logiskt
      1 logistiska
      1 logistiskt
      3 lögn
      1 lögnen
      3 lögner
      3 lögnerna
     12 logoped
      6 logopeden
      3 logopedens
      7 logopeder
      2 logopedexamen
      1 logopedförbundet
      2 logopedi
      5 logopedisk
      2 logopediska
      1 logopediskt
      2 logopedutbildning
      1 logopedutbildningen
      1 logopedyrket
      7 logos
      3 logotyp
      3 logotypen
      1 lohr
      1 lojala
      1 löjliga
      1 löjtnant
      1 löjtnantshjärta
      1 löjtnantshjärtesläktet
      6 lök
     50 lokal
     50 lokala
      2 lokalanestetika
      1 lokalbedövad
      1 lokalbedövar
     24 lokalbedövning
      1 lokalbedövningen
      2 lokalbedövningsmedel
      3 lokalbedövningsmedlet
      1 lokalbefolkning
      1 lokalbefolkningen
      1 lokalbehandla
      6 lokalbehandling
      1 lokalen
     14 lokaler
      2 lokalerna
     11 lokalisation
      3 lokalisationer
      7 lokalisera
     16 lokaliserad
      4 lokaliserade
      1 lokaliserades
      2 lokaliserar
      2 lokaliseras
      5 lokaliserat
      2 lokalisering
      1 lokaliseringsmärken
      1 lokalreaktioner
      1 lokalrengöring
     35 lokalt
      1 lokaltiden
      3 lokalvård
      7 lokalvårdare
      2 lokalverkande
      3 lokan
      1 loke
      2 löken
      1 loket
      1 loketrätan
      1 lokförare
      1 löklik
      1 lokomotiv
      1 lokomotorisk
      1 lokor
      1 lökväxt
      3 lökväxter
      1 lolo
      1 lomanus
      1 lomb
      1 lomma
      3 lömsk
      1 lömska
      1 [l�on]
      2 lön
      1 lönar
     26 london
      1 londonpapyrusen
      1 londons
      1 lönearbete
      1 lönen
      1 löner
      5 long
      1 longipes
      1 longitudinal
      1 longitudinala
      2 longitudinalis
      2 longitudinell
      3 longitudinella
      1 löning
      1 lönn
      2 lönsamt
      2 lönskaläge
      2 look
      2 loop
      1 loopar
      1 loopdiuretika
      1 loopen
      1 loopformade
      1 loopileostomi
      2 loopmetoden
      1 löp
      3 löpa
      5 löpande
      1 löparbanor
      4 löpare
      1 löpares
      3 löparknä
      1 löpe
     45 löper
      1 loperamid
      1 lopid
     10 löpning
      1 löpningen
      5 lopp
      6 loppan
      1 loppans
      8 loppet
      9 loppor
      4 lopporna
      1 loppornas
      1 löpsteget
      2 löpt
      2 löpte
      1 löptid
      1 loquax
      1 lord
      1 lördagsgodis
      3 lordos
      1 lordosis
      1 lordotisk
      2 loreal
      1 lorenzo
      4 lorenzos
      1 lori
      1 lornjett
      5 los
     11 lös
     29 lösa
      1 lösandet
      3 lösare
      8 lösas
      1 lose
      1 losec
     24 löser
     20 löses
      1 lösgjorde
      1 lösgör
      1 lösgöras
      2 lösgörs
      3 löslig
      4 lösliga
      6 löslighet
      1 lösligheten
      8 lösligt
     49 lösning
     23 lösningar
      1 lösningarna
      1 lösningars
     20 lösningen
      1 lösnings
      1 lösningsförslag
     24 lösningsmedel
      1 lösningsmedelsångor
      1 lösningsmedelsorsakad
      1 lösningsmedlen
      2 lösningsmedlet
      1 lösögonfransar
      1 lösöret
     14 loss
      8 löss
      2 lossa
      1 lossade
      1 lossades
      2 lossar
      1 lossas
      1 lossat
      1 lössen
      4 lossna
      1 lossnade
     13 lossnar
      2 lossnat
      1 lost
     20 löst
      5 lösta
      1 löstagbar
      1 löstagbara
      1 löstagbart
      2 löste
      1 lösts
      6 lotion
      2 lotioner
      1 lotions
      1 lottades
      1 lottats
      2 loudness
     10 louis
      2 louise
      1 louisencefalitvirus
      1 louisiana
      1 loup
      1 loupgarou
      2 loups
      1 louyse
      2 lov
      6 löv
      6 lovande
      2 lovar
      1 lovärt
      1 love
      1 lovely
      3 löven
      2 lovestruck
      4 lövfällande
      1 lovis
      1 lövkojor
      1 lovligt
      1 lovordat
      1 lovplikt
      4 lövskog
      1 lövskogar
      1 lövskogs
      1 lövskogshällar
      1 lövskogsmarker
      1 lövskogsnunnan
      3 lövträd
      1 lovvärda
      7 low
      1 löwenhjelm
      1 lower
      1 löylyä
      1 loz�re
      4 lp
      2 lps
      1 lqts
      1 lrv
     33 lsd
      1 lsdbruk
      1 lsdpåverkan
      1 lsdrus
      1 lsdterapi
      1 lsdupplevelsen
      1 lsekretet
      5 lss
      1 lsystemet
      1 lta
      1 ltp
      1 lubowe
      6 lubrikation
      6 lubrikationen
      1 lubrikerade
      1 lubuko
      1 lubulära
      3 luc
      1 lucid
      4 lucka
      1 luckan
      2 luckor
      1 luckra
      1 ludd
      1 ludda
      1 luddiga
      1 luden
      4 ludvig
      3 ludwig
      1 ludwigsburg
      1 ludwigshafenoppau
      1 luecke
      1 lues
    107 luft
      1 lufta
      1 luftbeständiga
      1 luftbh
      1 luftblandning
      1 luftblåsa
      1 luftblåsor
      1 luftbubbla
      1 luftbubblor
      3 luftburen
      2 luftburet
      8 luftburna
      1 luftdriven
      3 luftemboli
      1 luftembolier
     55 luften
      7 luftens
      1 lufterian
      1 lufterianer
      1 lufterianerna
      1 luftfarkoster
      3 luftflöde
      4 luftflödet
      1 luftföreningar
      1 luftförorening
      7 luftföroreningar
      2 luftfuktare
      8 luftfuktighet
      4 luftfuktigheten
      1 luftfylls
      1 lufthalter
      2 luftigt
      1 luftkanalerna
      1 luftkonditionering
      1 luftkonditioneringssystemet
      2 luftkuddar
      1 luftlandsattes
      1 luftmolekyler
      1 luftmotståndet
      1 luftningen
      2 luftningsbassängen
      1 luftningsbassänger
      1 luftningsbassängerna
      1 luftombyte
      1 luftomsättningen
      1 luftpassage
      2 luftpassagen
      1 luftrenande
      9 luftrenare
      2 luftrenaren
      6 luftrening
      1 luftreningen
      3 luftrör
      8 luftrören
      2 luftrörens
      1 luftröret
      1 luftrörsastma
      1 luftrörsbesvären
      1 luftrörskatarr
      1 luftrörsproblem
      1 luftrörsslemhinnan
      1 luftsäckarna
      2 luftslang
      1 luftslangen
      1 luftstöt
      2 luftströmmen
      2 luftstrupe
     26 luftstrupen
      3 luftstrupens
      2 lufttätt
      1 lufttemperaturen
      1 lufttomma
      2 lufttryck
      4 lufttrycket
      5 luftväg
     14 luftvägar
     75 luftvägarna
      6 luftvägarnas
      1 luftvågen
      2 luftvägen
      1 luftvägsavstängning
      1 luftvägsbesvär
      1 luftvägsepitel
      2 luftvägsepitelet
      1 luftvägshantering
      1 luftvägsinfekterade
      2 luftvägsinfektion
      9 luftvägsinfektioner
      2 luftvägsobstruktion
      1 luftvägsreaktioner
      2 luftvägssekret
      1 luftvägssjukdom
      1 luftvägssjukdomar
      1 luftvägsskydd
      1 luftvibrationer
      1 luftvolym
      1 luftvolymen
     13 lugn
      5 lugna
     28 lugnande
      1 lugnare
      5 lugnt
      1 luigi
      1 luk
      1 lukas
      1 lukes
      1 lukrativ
      1 lukrativa
     50 lukt
     10 lukta
      1 luktade
      1 luktämne
      1 luktämnen
      1 luktande
      5 luktar
      1 luktärt
      1 luktbanor
      1 luktblindhet
      1 luktbulben
      5 lukten
      1 luktepitelet
      5 lukter
      1 lukterna
      1 luktförmågan
      2 luktfri
      1 luktfria
      1 luktkänsliga
      3 luktlös
      1 luktlösa
      1 luktnerven
      1 luktproblem
      1 luktproblemen
      1 luktprov
      1 luktreducering
      2 luktsalt
      4 luktsinne
      6 luktsinnet
      1 luktstimuli
      2 lumbago
      1 lumbal
      1 lumbaldrän
     11 lumbalpunktion
      2 lumbalpunktionen
      2 lumbricoides
      6 lumen
      1 lumenala
      1 lumene
      1 lummerväxter
      1 lumpektomi
      1 lumpektomiingreppet
      1 lumpektomin
      1 lumps
      1 lunardo
     18 lund
      2 lundar
      1 lundbeck
      1 lundberg
      3 lundborg
      1 lundens
      1 lundin
      2 lundkvist
      6 lunds
      1 lundstr
      2 lundväxt
      1 lundväxter
      1 lunetiers
      2 lung
      8 lunga
      3 lungabscess
      2 lungabscesser
      1 lungadenocarcinom
     31 lungan
      5 lungans
      1 lungartären
      1 lungartärer
      1 lungbaserna
      6 lungblåsorna
      1 lungbristningar
     55 lungcancer
      1 lungcancer[]
      1 lungcancerfall
      1 lungcancerrisken
      2 lungcancersjukdomar
      1 lungcancertalk
      1 lungcancertumörer
      1 lungcancerutveckling
      2 lungcancrar
      6 lungcarcinom
      1 lungcirkulationen
      1 lungdel
     20 lungemboli
      1 lungembolier
      1 lungemfysem
      3 lungfibros
      1 lungförändringar
      1 lungfriska
      5 lungfunktion
      3 lungfunktionen
      5 lungfunktionsnedsättning
      2 lungfunktionsundersökning
      1 lunghjärtsjukdom
      1 lunginfiltrat
     90 lunginflammation
      4 lunginflammationen
      2 lunginflammationer
      1 lunginflammationsfallen
      2 lungkapacitet
      1 lungkapillärerna
      1 lungkärlens
      4 lungkollaps
      1 lungkomplikationer
      5 lungkretsloppet
      1 lungläkare
      1 lungläkaren
      1 lunglob
      3 lungloben
      1 lunglober
      1 lungmaskiner
      1 lungmognad
      2 lungmognaden
     12 lungödem
     28 lungor
    153 lungorna
     15 lungornas
      1 lungparenkymet
      2 lungpåverkan
      9 lungpest
      2 lungproblem
      1 lungpunktering
      4 lungräddning
     13 lungröntgen
     12 lungsäcken
      3 lungsäckens
      1 lungsäcks
      1 lungsäcksblad
      1 lungsäcksbladet
      1 lungsäcksförtjockning
      1 lungsäcksvävnad
     11 lungsjukdom
     14 lungsjukdomar
      1 lungsjukdomarna
      1 lungsjukdomcopd
      1 lungsjukes
      1 lungsjukgymnastik
      1 lungskada
      4 lungskintigrafi
      1 lungsot
      1 lungsprängning
      1 lungstrukturer
      1 lungtrakten
      6 lungtuberkulos
      1 lungtumör
      5 lungvävnad
      8 lungvävnaden
      1 lungvener
      4 lungvolym
      1 lungvolymen
      1 lunsford
      1 lunta
      1 luntlapp
      3 lupus
      2 lura
      1 lurar
      1 lurarna
      1 luras
      1 lurat
      1 lurias
      1 lusbräda
      2 lusbrädan
      2 lusen
      2 lusflugor
     14 lust
      1 lustan
      2 lustar
      4 lusten
      1 lustfyllda
     22 lustgas
      3 lustgasen
      1 lustgasrus
      1 lustgassystem
      1 lustprincipen
      1 lustsjukan
      1 lustupplevelserna
      1 luta
      1 lutad
      2 lutande
      8 lutar
      9 luteiniserande
      1 luteiniseringhormon
      1 luteom
      1 lutetia
      1 luteum
      1 luteus
      1 luther
      1 luthersk
      1 lutherska
      3 lutning
      1 lutningar
      1 lutningen
      1 lutningsförändring
      1 lutstänk
      1 lutsträngar
      1 lützenberg
      2 lux
      4 luxemburg
      1 luxuöst
      1 lv
      1 lvfs
      1 l�v�ya
      1 lycicus
      8 lycka
      7 lyckad
     11 lyckade
     35 lyckades
     25 lyckas
      1 lyckat
     30 lyckats
      1 lycklig
      2 lyckligare
      1 lyckligt
      5 lyckligtvis
      1 lyckoamuletter
      1 lyckobringande
      2 lyckosam
      1 lyckosamt
      1 lyckosubstanser
      2 lycoctonum
      1 lycosa
      1 lyda
      1 lydde
      6 lyder
      1 lydisk
      1 lydiske
     12 lyft
      7 lyfta
      1 lyftarmuskel
      2 lyftas
      4 lyfte
     19 lyfter
      4 lyfts
      1 lyftselar
      1 lyftsele
      1 lyftsituationer
      1 lyhörda
      1 lyhördhet
      3 lykopen
      1 lyktstolpe
      5 lyme
      1 lymecyklin
      3 lymerix
      2 lymfa
      2 lymfan
      1 lymfangiom
      1 lymfangiomgenetisk
      1 lymfangiosarkom
      8 lymfatisk
      8 lymfatiska
      2 lymfatiskt
      1 lymfbanorna
      7 lymfkärl
      3 lymfkärlen
      1 lymfkärlssystemet
      1 lymfknuta
      9 lymfknutor
      2 lymfknutorna
      1 lymfkörtelförändringar
      1 lymfkörteln
     10 lymfkörtlar
      6 lymfkörtlarna
      1 lymfkörtlarskelett
      1 lymfnoder
      1 lymfnoderna
      1 lymfnodscancer
      1 lymfoblastisk
      2 lymfocyt
      1 lymfocytär
      1 lymfocyten
     14 lymfocyter
      4 lymfocyterna
      2 lymfocytisk
      3 lymfödem
      1 lymfografi
      1 lymfoid
     27 lymfom
      2 lymfomen
      1 lymfomprognosen
      1 lymfoplasmocytiskt
      4 lymfsystemet
      2 lymfvätska
      1 lymfvätskan
      3 lymfvävnad
      1 lymfvävnaden
      2 lymphadenopathyassociated
      1 lymphoma
      1 lynnet
      1 lynnighet
      1 lyomyces
      2 lyon
      5 lypsyl
      1 lyrica
      2 lyrisk
      1 lys
      2 lysa
      2 lysande
      1 lysatreaktioner
      1 lysdioder
      2 lyser
      2 lyserar
      1 lyseras
      1 lysergsäurediethylamid
      2 lysergsyra
      3 lysergsyradietylamid
      1 lysholm
      3 lysin
      1 lysis
      1 lysosom
      1 lysrör
      1 lyssa
      1 lyssavirus
     11 lyssna
      2 lyssnade
      1 lyssnades
      1 lyssnande
      1 lyssnandet
      3 lyssnar
      3 lyssnare
      1 lyssnarna
      1 lyssning
      3 lyssningshjälpmedel
      1 lysten
      1 lysved
      1 lyx
      1 lyxiga
      1 lyxzén
     86 m
      4 �m
      3 ma
     16 må
      1 maa
      1 määttä
      4 mabthera
      2 mabuse
      2 mac
      1 macadamianötter
      2 macchiarelli
      1 macdonald
      1 macdonaldtriaden
      1 macfarlan
      1 machine
      1 machupo
      1 macintoshblad
      1 macleod
      1 macrolepiota
      1 macropinocytos
      1 macropus
      1 macrostachys
      1 macula
      1 maculans
      1 macvärdet
      1 mad
      2 madagaskar
      1 madams
      2 madeira
      1 madeiraflädern
      1 madhava
      1 madness
      1 madnessång
      3 madonna
      1 madrasser
      2 madrid
     22 mag
      1 magåkomma
      2 magasin
      2 magazine
      5 magbesvär
      2 magbiverkningar
      1 magbråck
      2 magcancer
      3 magdelarna
     16 mage
      1 magement
     43 magen
      5 magens
      1 mager
      1 magerhet
      1 magert
      1 maggie
      1 maggropen
      6 magi
      3 magic
      1 magiker
      1 magikers
      1 maginfektion
      1 maginfluensa
      3 maginnehåll
      5 maginnehållet
      1 maginnehållets
      1 magisk
     13 magiska
      1 magiskreligiösa
      5 magiskt
      2 magister
      3 magisterexamen
      2 magkatarr
      1 magkatarrliknande
      1 magknip
      1 magkramp
      1 magkramper
      3 magmatiska
      7 magmunnen
      1 magmuskel
      1 magnavox
      4 magnecyl
     13 magnesium
      1 magnesiumammoniumfosfat
      2 magnesiumbrist
      1 magnesiumjon
      1 magnesiumjoner
      1 magnesiumoxid
      1 magnesiumrik
      1 magnesiumrika
      1 magnesiumsalter
      1 magnesiumsilikatklorit
      1 magnesiumstearat
      1 magnesiumsulfat
      2 magnesiumvärdena
      1 magneter
      1 magnetfält
      7 magnetisk
      6 magnetiska
      1 magnetiskt
      3 magnetism
      6 magnetkamera
      1 magnetkameraangiografi
      4 magnetkameraundersökning
      1 magnetresonans
      9 magnetresonanstomografi
      1 magnetröntgen
      1 magnonmänniskan
      5 magnus
      1 magnusekenenstierna
      1 magoch
      7 magont
      1 magoperationer
      6 magproblem
      1 magproblemen
      1 magpumpning
      1 magra
      1 magraste
      3 magsäck
     80 magsäcken
      5 magsäckens
      1 magsäcks
      8 magsäckscancer
      1 magsäcksinflammation
      1 magsäckskroppen
      1 magsäcksslemhinnan
      3 magsaft
      2 magsaften
     10 magsår
      1 magsåret
      1 magsårssjukdomar
     11 magsjuka
      1 magsjukan
      1 magsjukdom
      1 magsjukesymtom
      6 magsmärta
      9 magsmärtor
      3 magstärkande
      1 magstrupe
      1 magstrupen
      4 magsyra
      1 magsyran
      1 magsyrans
      1 magsyretåligt
      1 magtarmbesvär
      1 magtarminflammationer
      2 magtarmkanal
      1 mag�tarmkanal
     20 magtarmkanalen
      1 magtarmkanalens
      1 magtarmkatarr
      1 magtarmsjukdom
      1 magtarmsystemet
      1 magtömning
      1 magtrakten
      2 magvärk
      1 mahabharata
      3 måhända
      1 maharishi
      1 maharishis
      1 mahesh
      1 mahler
      3 maiden
      1 maidenform
      2 maieutik
      1 maile
      1 maillardreaktionen
      1 maimonides
      2 main
      1 mainstream
      1 mainstreamkultur
      1 mainstreamkulturen
      1 mainstreampsykiatrin
      1 maintainability
      2 maintenance
      2 maintenaz
      5 maitenaz
     30 maj
      2 majalis
      1 majevtik
      1 majja
      1 majjuni
      3 majonnäs
      5 major
     11 majoritet
     26 majoriteten
      1 majoritetsbefolkningen
     10 majs
      1 majsen
      1 majsolja
      1 majspåsar
      3 majsstärkelse
      1 majsstärkelsepuder
      1 majsvälling
      2 majus
      1 mak
      1 makabra
      1 makalös
      1 makarmakor
      1 makarnas
      1 make
      1 makedonien
      6 maken
      2 makeup
      1 makeupartister
      1 makololofolket
      1 makroadenom
      1 makrobiotik
      1 makrobiotiken
      1 makrocyterna
      1 makrofag
      2 makrofagen
     19 makrofager
      2 makrofagerna
      1 makrofagernas
      1 makrogametofyten
      1 makrogamofyten
      2 makroglobulinemi
      1 makrokosmos
      1 makrolid
      7 makrolider
      1 makromolekylära
      1 makromolekylärt
      2 makromolekyler
      3 makronutrienter
      1 makros
     15 makt
      1 mäktar
      3 makten
      3 makter
      1 makters
      1 maktfaktor
      1 mäktig
      1 mäktiga
      1 mäktigaste
      1 maktinstrument
      2 maktlöshet
      1 maktlöst
      1 maktmedel
      1 maktobalansen
      1 maktposition
      1 maktutövning
      3 makula
      1 makulopapulösa
      5 mal
     67 mål
      1 mala
      1 måla
      7 malabsorption
      1 malabsorptionssjukdomar
      1 målad
      1 maladaption
      2 maladaptiva
      6 målade
      1 malajer
      2 malajerna
      2 malajiska
      1 malandanti
      2 målande
      1 malar
      3 målar
      1 målare
      1 målaren
      1 mälaren
      4 målarfärg
      1 målarfärgen
     48 malaria
      2 malariacykeln
      1 malariadrabbade
      1 malariadrabbat
      1 malariae
      1 malariainfektion
      1 malariamedel
      1 malariamedicin
      1 malariamyggan
      1 malariamyggor
      1 malariamyggorna
      3 malarian
      1 malariaparasiten
      2 malariaparasiter
      1 malariasmittan
      1 malariaspridande
      1 malariasymptomen
      2 malariatillfällen
      1 malarone
      1 mälartrakterna
      2 målas
      4 målat
      1 malawi
      2 malayi
      1 malaysia
      1 malberg
      1 målbeskrivningen
      1 målbrott
     14 målbrottet
      2 målbrottsstörning
      1 målcellen
      6 målceller
      3 målcellerna
      1 malcolm
      1 mald
      1 malda
      1 malde
      1 maldescenderade
      2 maldi
      1 maldigestion
      1 male
      6 målen
      1 måleri
     23 målet
      1 måletmålen
      1 målets
      1 malformation
      1 målgrupp
      1 målgrupper
      1 malheim
      1 malheims
      1 malheur
      3 mali
     24 malign
     18 maligna
      2 malignitet
      2 maligniteter
      5 malignt
      1 målinriktade
      1 målinriktat
      1 malkulor
      2 mall
      1 mallei
      1 malleus
      4 mallophaga
      1 mallophagerna
      1 mallorca
      1 malmedel
      2 målmedveten
      1 malmen
      2 malmer
     14 malmö
      1 målmolekylen
      3 målning
      3 målningar
      1 målningarna
      1 målningsarbeten
      2 malnutrition
      1 malocklusioner
      2 målområdet
      2 målorgan
      1 målorganet
      1 malört
      1 malpighiska
      3 mals
      2 målsättning
      5 målsättningar
      5 målsättningen
      1 målskytte
      5 malt
      3 malta
      1 maltamylaserna
      1 måltavla
      1 måltavlor
      1 maltextrakt
      1 malthus
     16 måltid
      4 måltiden
      1 måltidens
     12 måltider
      2 måltiderna
      1 måltidsobservation
      1 mältningen
      4 maltos
      1 maltoscannabis
      1 malttorka
      1 måltumören
      1 måltumörens
      1 målvävnad
      1 målvävnader
      1 målvävnaderna
      2 målvikt
      1 målyta
      1 malzieu
      1 mamba
      1 mameluckerna
      1 mamillosa
      1 mamma
      1 mammae
      1 mammakläder
      8 mamman
      2 mammans
      1 mammografer
     16 mammografi
      1 mammogram
      1 mammogrammet
      1 mammor
      1 mammorna
      1 mammosite
      1 mammoth
      1 mamsa
   3381 man
     31 mån
    392 män
     10 mana
      1 måna
     30 månad
      7 månaden
    161 månader
     10 månaderna
     18 månaders
      2 månadersperiod
      1 månadsgammalt
      1 månadskopp
      1 månadslånga
      1 månadslinser
      4 management
      1 månar
      2 månatlig
      1 månatligt
      1 manchester
      1 manchuerna
      1 mandat
      2 mandel
      1 mandelmjölk
      1 mandibelframdragande
      1 mandibular
      2 mandlar
      2 mandragora
      1 mandragoraroten
      3 månen
      3 manet
      4 maneten
      1 manetens
      7 maneter
      1 manetliknande
      1 maneuver
      1 manev
      1 manfred
      1 mang
      4 manga
   1039 många
      2 mangan
      2 mangandioxid
      1 manganviioxid
      1 mångårig
      1 mångårigt
      1 mångas
    164 mängd
     99 mängden
      1 mångder
    127 mängder
      1 mängderna
      1 mångdimensionell
      1 mångdimensionella
      2 mångdubbelt
      1 mångdubblas
      1 mangeais
      2 mangel
      1 mangelbodar
      1 mangelbräde
      2 mangelbräden
      1 mängen
      1 mangeons
      1 manger
      3 mångfald
      2 mångfalden
      1 mångfaldigar
      2 mångformig
      1 mångfröig
      1 mangling
      1 mångmiljonbelopp
      3 mango
      1 mångsidig
      2 mångt
      3 mångtydig
      1 mångtydiga
      1 mångtydigt
      3 manhattan
      1 manhunters
     17 mani
      3 mania
      6 manier
      1 manifest
      1 manifesta
      1 manifestation
      3 manifestationen
      4 manifestationer
      1 manifesterade
      6 manifesterar
      5 manifesteras
      2 manifesterat
      6 manikyr
      1 manikyrbehandlingar
      1 manin
      5 maniok
      1 maniokberedningen
      1 maniokmjöl
      1 maniokodlande
      1 maniokrötter
      1 manioksorter
      7 manipulation
      1 manipulationens
      2 manipulativ
      1 manipulativa
      1 manipulative
      1 manipulativt
      5 manipulera
      1 manipulerade
      1 manipulerandet
      1 manipulerar
      2 manipuleras
      2 manipulerat
      1 manipulering
      1 manipulus
      3 manisk
      1 maniska
      1 manitoba
      1 mänkvinnor
     25 manlig
     44 manliga
     15 manligt
      1 manligtvuxet
      1 manna
      1 mannans
      1 mannekänger
     36 mannen
     18 männen
      2 mannenpojken
     15 mannens
      3 männens
    134 människa
      1 människamaskinsystem
    191 människan
     95 människans
     19 människas
      2 människo
      1 människoapor
      1 människoaporna
      1 människoapornas
      1 människoblod
      1 människoceller
      1 människoföda
      1 människohår
      1 människohjärtats
      1 människohuvud
      3 människokropp
      3 människokroppar
     24 människokroppen
      6 människokroppens
      1 människokunskap
      2 människoliv
      1 människoloppan
      1 människooffer
      2 människoorsakade
    728 människor
      1 människoraser
      1 människorättskämpen
      8 människorna
      2 människornas
      1 människorref
     39 människors
      1 människosjälen
      1 människoskapat
      3 människosläktet
      1 människosläktets
      1 människospermien
      2 människosyn
      1 människovärdiga
      1 mannitol
      1 mannos
      3 manodepressiv
      3 manodepressivitet
      1 manometer
      1 manövern
      1 manöverpanel
      1 manövrera
      1 manövrerar
      1 manövreras
      5 mans
      2 måns
      7 mäns
      1 mansfield
     27 mänsklig
     54 mänskliga
      6 mänskligheten
      2 mänsklighetens
     11 mänskligt
      1 manskön
      2 mansonia
      1 mantakassa
      1 mantalsskriven
      1 mantegazza
      3 mantegazzianum
      2 mantel
      1 manteldjuren
      1 mantimme
      1 mantoux
      1 mantouxtest
      4 mantouxtestet
      1 mantra
      3 mantran
     13 manual
      1 manualbaserad
      1 manualbaserade
      1 manualbaserat
      3 manualen
      4 manualer
      1 manuel
     11 manuell
      7 manuella
     11 manuellt
      1 manus
      1 manutergium
      2 mao
      2 maobhämmaren
      1 map
      1 mapkerksignaltransduktionsvägen
      1 maple
      1 maquet
     13 mår
      1 mara
      2 maran
      1 marantz
      1 marasm
      1 marasmer
      1 marasmiaceae
      1 marburg
      4 marburgvirus
      3 marcel
      1 marco
      1 marcus
      1 mårdhund
      4 mardröm
      5 mardrömmar
      4 maréchaussée
      1 maréchaux
      1 mareridt
      1 mareritt
      2 marfans
      2 märg
      1 marga
      4 margaret
      1 margareth
      3 margarin
      2 margarine
      1 margarinet
      1 margarinföretaget
      1 margarinproducenten
      1 märgel
      1 märgelsten
     16 märgen
      1 märgens
      1 märghålan
      3 marginal
      1 marginaleslentiformesbr
      1 marginaliserade
      1 marginalisering
      2 marginalområdet
      4 marginell
      3 marginellt
      2 margit
      1 margot
      1 märgspik
      6 maria
      1 marianne
      1 mariano
      6 marie
      1 marieberg
      1 mariestad
      1 marin
      2 marina
      1 marinakustik
      1 marinbiologi
      1 marinläkaren
      1 marinor
      1 marinpolisen
      1 marint
      1 marinum
      1 marion
      1 maritime
      2 maritimus
     22 mark
      5 märka
     16 markant
      1 markanta
      4 märkas
      8 märkbar
      2 märkbara
      4 märkbart
      1 markburen
     14 märke
     28 marken
      9 märken
      3 märkena
      3 marker
     16 märker
      4 markera
      2 markerad
      5 markerade
      2 markerar
      2 markeras
      1 markerat
      2 markeringar
      1 markerna
      1 märkesflikar
      1 märkesmedvetenheten
      1 märkesnamn
     11 märket
      1 markförstöring
      1 markledningar
      1 marklevande
      2 märklig
      3 märkliga
      2 märkligt
      2 marknad
     49 marknaden
      1 marknader
      1 marknadsanalys
      1 marknadsbolag
      1 marknadsför
      3 marknadsföra
      2 marknadsföras
      2 marknadsförde
      6 marknadsfördes
      9 marknadsföring
      2 marknadsföringen
      1 marknadsföringstillståndet
      6 marknadsförs
      1 marknadshandel
      1 marknadsledande
      1 marknadsundersökningar
      1 marknatsföring
      6 märkning
      1 märkningar
      4 märkningen
      1 marknivå
      1 markoch
     11 markör
      2 markören
      3 markörer
      2 markörerna
      1 markovkohortmodell
      1 markradonhalten
     18 märks
      1 märksamma
      3 märkt
      7 märkta
      1 marktäckare
      4 märkte
      2 märktes
      1 märkts
      1 marktschreyeri
      1 märkvärdiga
      1 märkvärt
      1 markytan
      1 marlboros
      1 marlene
      1 marlon
      1 marmor
      1 marmoratus
      2 marmorerad
      1 marmoreringar
      1 marmorskivor
      1 marocko
     29 mars
      1 marschera
      1 marscherade
      1 marseille
      1 marseilletvål
      1 marsh
      1 marshskalan
      2 marsilio
      1 marskalkämbetets
      3 marsvin
     12 martin
      1 martinieffekten
      1 martröð
      2 martyrskap
      1 marx
      1 marxistisk
      7 mary
      2 maryland
      1 masada
      3 mascara
      1 mascaran
     13 mask
      2 maskägg
      1 maskangrepp
      9 maskar
      8 maskarna
      4 maskarnas
      1 maskartade
      1 maskarter
     20 masken
      1 maskera
      1 maskerad
      1 maskerader
      1 maskerna
      3 maskformiga
      2 maskformigt
     10 maskin
      2 maskindisk
      1 maskinell
     17 maskinen
      2 maskinens
     13 maskiner
      1 maskineri
      1 maskinerna
      1 maskininstallationer
      1 maskinläsbar
      1 maskinrullning
      1 maskinskrivning
      1 maskmaterial
      1 maskopi
      1 masksjukdom
      1 maskulinisation
      1 maskulinitet
      1 masmovägen
      1 masochism
      2 mass
     20 massa
      3 massachusetts
      2 massäck
     23 massage
      1 massagebänk
      1 massagebehandlingar
      6 massagen
      1 massagens
      1 massageolja
      1 massagetekniker
      2 massaindustrin
      1 massajerna
      2 massakern
      1 massaladdning
      3 massan
      2 mässan
      1 massanalysator
      1 massanalysatorer
      1 masséin
      1 massenhet
      4 massera
      1 masserade
      2 masseras
      1 masseter
      1 massförgiftningar
      2 massgrav
      3 mässing
      7 massiv
      2 massiva
      2 massivt
      1 massladdning
      2 massladdningsförhållande
     38 mässling
      2 mässlingen
      1 mässlingens
      1 mässlings
      1 mässlingsepidemi
      1 mässlingsepidemier
      1 mässlingsfall
      1 mässlingsförekomsten
      1 mässlingsliknande
      1 mässlingspatienter
      1 mässlingsstammar
      8 mässlingsutbrott
      1 mässlingsvaccin
      1 mässlingsvaccination
      1 mässlingsvaccinet
      1 mässlingsvirus
      2 mässlingsviruset
      1 mässlingsvirusinfektion
      1 mässlingvirus
      1 mässlingviruset
      3 massmedia
      1 massmedial
      1 massmediebilder
      2 massmedier
      2 massmord
      4 massor
      1 massoterapi
      1 massövervakning
      1 massövervakningssamhälle
      2 masspektrometrar
      2 masspektrometri
      1 masspektrum
      1 massproducera
      1 massproducerade
      1 massproducerades
      1 massproduceras
      2 massproduktion
      2 masspsykos
      2 masstillverka
      1 masstillverkade
      1 masstillverkas
      1 massvaccination
      1 massvaccinering
      1 massvält
      3 mästare
      1 mästarnas
      1 mastcell
     12 mastceller
      2 mastcellerna
      2 mastcellsdegranulering
    335 måste
      7 mastektomi
      5 master
      1 mäster
      3 masterexamen
      1 masterprogrammet
      1 masters
      1 mastersexamen
      1 mastersutbildningar
      1 masterutbildningar
      3 mastit
      2 mastocytos
      1 mastodeton
      6 mastodyni
      4 mastoidit
      6 mastomys
      1 mastos
      5 masturbation
      1 masurien
      1 masurium
    139 mat
      1 mata
     88 mäta
      1 matade
      1 matades
      2 mataffärer
      1 matallergier
      1 matallergieri
      1 matar
      2 mätare
      3 mätaren
      1 mätarfabrikör
      2 matas
     32 mätas
      1 mätbar
      7 mätbara
      2 mätbart
      1 matberedning
      1 matberedningsytorna
      1 matbestick
      1 matbeteende
      1 matbistånd
      1 matbitar
      1 matbordet
      2 matbrist
      3 match
      1 matcha
      3 matchande
      2 matchar
      1 matchas
      1 matchat
      2 mätdata
      1 mätdon
      2 mate
      1 maté
      1 matein
      8 matematik
      1 matematikern
      1 matematikfärdigheter
      1 matematikprov
      2 matematiksvårigheter
      3 matematisk
      4 matematiska
      1 matematiskstatistisk
      3 matematiskt
     49 maten
      2 matens
      1 mater
     58 mäter
      4 materia
    128 material
      1 materialen
     39 materialet
      2 materialets
      1 materialism
      1 materialnamnet
      1 materialprov
      1 materialprovning
      1 materials
      1 materialt
      1 materialtjocklek
      1 materialvetenskap
      1 materias
      3 materiel
      2 materiell
      6 materiella
      1 materien
      1 materier
      1 mätfallanvändningsområden
      2 matfett
     20 matförgiftning
      1 matförgiftningar
      2 mathållning
      1 mathé
      1 mathew
      1 mathisen
      1 matindustrin
     11 mätinstrument
      2 matintag
      1 matintaget
      1 matkoma
      1 mätkretsar
      1 matkulturer
     14 matlagning
      3 matlagningen
      1 matlagningsgrädde
      1 matlagningshygien
      1 matlagningsmetod
      1 matlagningsmetoder
      1 matleda
      1 matledaillamående
      1 matledskvistar
      1 matluktsmak
      2 matlust
      1 matmärken
      4 mätmetod
      3 mätmetoder
      1 matnedbrytningen
     33 mätning
     28 mätningar
      2 mätningarna
      8 mätningen
      1 mätnoggrannheten
      1 matolja
      6 mätområde
      1 mätområden
      1 mätområderna
      1 matpartiklar
      1 matporslin
      2 maträtter
      7 matrester
      1 mätresultaten
      2 matris
      1 matriser
      5 matrix
      1 matrixet
      1 matrixmetalloproteaser
      3 mats
     33 mäts
      2 matsäck
      1 matsäkerheten
      1 matsäkerhetsmyndighet
      1 mätsignal
      2 mätsignalen
      1 matskedar
      3 matsmältning
      6 matsmältningen
      1 matsmältnings
      2 matsmältningsenzymer
      1 matsmältningsfaser
      2 matsmältningskanal
     10 matsmältningskanalen
      1 matsmältningskanalens
      2 matsmältningsprocessen
      2 matsmältningssystem
      3 matsmältningssystemet
      3 matspjälkning
      4 matspjälkningen
      1 matspjälkningsenzymer
      1 matspjälkningskanal
      1 matspjälkningskanalen
      2 matspjälkningssystem
      3 matspjälkningssystemet
      1 matstationer
      1 mätstörningar
      4 matstrupe
     47 matstrupen
      1 matstrupens
      3 matstrupscancer
      1 matstrupsmunnenesofagussfinktern
      7 matsvamp
      1 matsvampar
      4 matt
     46 mått
      8 mätt
      3 matta
      1 mättad
      2 mättade
      1 måttagning
      2 mattas
      1 mättas
     12 mättat
      1 mattats
      1 matte
      1 mätte
      2 mättekniker
      7 måtten
      1 måttenheten
      6 måttet
      2 matteusevangeliet
      1 måttfulla
      1 måttfullhet
      2 matthet
      2 matthew
      2 matthias
      1 matthiesen
      1 mättid
     27 måttlig
      7 måttliga
      1 måttlighet
      2 måttligt
      1 måttmässigt
      4 mättnad
      1 mättnadsdykning
      1 mättnadsgrad
      1 mättnadshormon
      1 mättnadskänsla
      1 mättnadsreglerande
      1 måtto
      2 mattor
      1 måttstock
      1 måttsy
      1 måttsystemet
      1 mätuppgiften
      1 maturity
      1 mätutrustning
      1 matvägran
      1 matval
      7 matvanor
      1 matvanorna
      2 matvaran
      3 mätvärde
      6 mätvärden
      2 mätvärdet
     10 matvaror
      1 matvarorna
      1 maud
      2 maurice
      2 mauvein
     15 max
      1 maxfactor
      1 maxhastighet
      1 maxibindor
      1 maxillasis
     10 maximal
     10 maximala
      7 maximalt
      2 maximera
      1 maximerat
      2 maximum
      1 maximumintensity
      1 maxin
      1 maxpuls
      1 maxpulsen
      1 maxspänning
      1 may
      1 mayafolket
      4 mayaindianerna
      1 mayaperioden
      1 maybelline
      1 mayer
      1 mayerrokitanskyküsterhausersyndrom
      2 mazess
      2 mb
      2 mbd
      1 mbensendiol
      2 mbp
      1 mbsr
      1 mbt
      1 mccann
      1 mcclintockeffekten
      1 mcdowell
      1 mci
      2 mckenzie
      1 mcm
      1 mcpherron
      1 mcr
      1 mcv
      3 md
      1 mda
      1 mdihydroxibensen
      1 me
      1 meagans
      1 meal
      1 measles
      1 measurement
      1 meat
      2 mebendazol
      2 meca
      2 mecfs
      1 mecfspatienter
      1 mechanism
      1 mecka
      1 meckels
      1 meconopsis
   8488 med
      1 medaljen
      2 medaljer
    468 medan
      1 medans
      1 medantibiotikaresistensavses
     14 medarbetare
      1 medarbetares
      2 medarbetarna
      1 medarbeterska
     14 medborgare
      1 medborgarens
      2 medborgarna
      1 [medborgarnas]
      1 medborgarorganisationer
      1 medbrottsling
      3 meddela
      1 meddelande
      7 meddelanden
      2 meddelandena
      1 meddelandet
      1 meddelar
      1 meddelas
      3 meddelat
      2 médecine
    185 medel
      8 medelåldern
      7 medelålders
      2 medelartärtryck
      1 medelbentäthetsvärdet
      1 medelcellvolym
      1 medelengelska
      1 medelgod
      1 medelhalten
      6 medelhavet
      1 medelhavsdiet
      4 medelhavsdieten
      1 medelhavskost
      2 medelhavsländer
      6 medelhavsområdet
      1 medelhavsregionen
      1 medelhög
      1 medelhöga
      1 medelinkomstländer
      2 medelklassen
      1 medelklassfamiljer
      1 medelkoncentrationen
      3 medellängden
      1 medellångt
      2 medellinjesnitt
      8 medellivslängd
      1 medellivslängder
      1 medelljudnivån
      1 medelnivå
      2 medelpersonen
      1 medelpunkt
      1 medelresultat
      6 medelst
      1 medelstark
      1 medelstarka
      3 medelstora
      2 medelstort
      2 medelsvår
      1 medelsvåra
      3 medeltal
      3 medeltid
     10 medeltida
     32 medeltiden
     11 medeltidens
      1 medeltidsbaden
      2 medeltidslatin
      4 medelvärde
      1 medelvärden
      6 medelvärdet
      1 medelvarma
     40 medfödd
     43 medfödda
      4 medföljande
      1 medföljde
      1 medföljer
     87 medför
     38 medföra
      1 medförande
      1 medförare
      6 medförde
      1 medförfattare
      3 medfört
     17 medfött
      1 medgav
      1 medge
     10 medger
      1 medges
      1 medgett
      1 medgivet
      1 medha
      1 medhjälp
     27 media
      1 mediaflödet
      3 medial
      4 medialt
      1 mediana
      2 medianåldern
      1 medianinsatstiden
      2 medianöverlevnaden
      1 medianpris
      1 medianus
      2 medianusnerven
      1 mediastinala
      2 mediastinalemfysem
      1 mediastinalt
      3 mediastinum
      1 mediator
      6 mediatorer
      1 mediatorsubstanser
     19 medical
      1 médicale
      1 medicering
    147 medicin
      1 medicinala
      1 medicinalansvarskommitten
      1 medicinalförfattningar
      1 medicinalförfattningarna
      2 medicinalis
      1 medicinalkol
      1 medicinallag
      1 medicinallagar
      1 medicinalpersonal
      3 medicinalstyrelsen
      1 medicinalstyrelsens
      1 medicinalsystem
      5 medicinalväxt
      4 medicinalväxter
      1 medicinalväxters
      2 medicinare
      1 medicinaren
      1 medicinarkåren
      1 medicinartad
      1 medicinbibliotek
      2 medicinboll
      2 medicinbollar
      1 medicinbollen
      1 medicindrog
     13 medicine
     69 medicinen
      3 medicinens
     67 mediciner
      3 medicinera
      1 medicinerade
      3 medicineras
      1 medicinerat
      2 medicinerats
     57 medicinering
      2 medicineringar
      7 medicineringen
      9 medicinerna
      1 medicines
      1 medicinflaskor
      1 medicinförpackningar
      1 medicinfria
      1 medicinhistoria
      1 medicinhistorien
      1 medicinhistoriens
      1 medicinhistoriskt
      1 medicinman
      1 medicinmän
    221 medicinsk
    206 medicinska
      1 medicinskakliniska
     77 medicinskt
      1 medicinsktbiologiska
      1 medicinstudent
      2 medicinstudenter
      1 medicinteknisk
      4 medicintekniska
      1 medicintekniskt
      1 medicintidskriften
      1 medicintillfällen
      1 medicintillförsel
      2 medicinvetenskapen
      1 medicis
      6 medicum
      1 mediemogul
      8 medier
      4 medierar
      3 medieras
      1 mediers
      1 mediet
      1 medikalisering
      1 medimix
      1 medimmunhämmande
      2 medinensis
      1 medinska
      1 mediokra
     35 meditation
      2 meditationen
      2 meditationens
      1 meditationer
      1 meditationsformer
      2 meditationsmetod
      1 meditationsövningar
      1 meditationsposer
      1 meditera
      1 mediterar
      1 mediterranei
      1 mediterraniae
      8 medium
      1 medkännande
      9 medkänsla
      2 medlare
      6 medlem
     35 medlemmar
     11 medlemmarna
      1 medlemmen
      1 medlemsförbund
      2 medlemskap
      1 medlemskapet
      3 medlemsländer
      2 medlemsländerna
      1 medlemsländernas
      5 medlemsstater
      4 medlemsstaterna
      8 medlen
     33 medlet
      1 medlets
      1 medlidande
      3 medline
      2 medmänniska
      1 medmänniskor
      1 medräknade
      1 medströms
      1 medtunntarmensinnehåll
      6 medulla
      4 medullär
      1 medulloblastom
      2 medusa
      1 medusae
      1 medusans
      1 medusatyp
      3 medusor
      1 medvandrande
      6 medverka
      1 medverkan
      9 medverkar
     15 medvetande
      1 medvetandedjup
      1 medvetandeförlust
      1 medvetandeformer
      1 medvetandegör
      2 medvetandegöra
      7 medvetandegrad
      4 medvetandegraden
      1 medvetanden
      1 medvetandenivå
      2 medvetandepåverkan
      1 medvetanderubbning
      1 medvetanderubbningar
      2 medvetandesänkning
     14 medvetandet
     12 medvetandetillstånd
     32 medveten
      1 medvetendegrad
     10 medvetenhet
      3 medvetenheten
      1 medvetenhets
      1 medvetenhetsutvecklad
     12 medvetet
     18 medvetna
      7 medvetslös
      2 medvetslösa
     23 medvetslöshet
      1 medvetslöst
     12 mefedron
      1 megakaryocyt
      1 megapodiidae
      1 meget
      1 megmagnetoencephalography
      1 mehmet
      3 mei
      1 meiinnehållet
      1 meijer
      1 meijirestaurationen
      4 meios
      2 meiosen
      1 meioserna
      7 mejeriprodukter
      1 mejl
      1 mekanik
     18 mekanisk
     16 mekaniska
     18 mekaniskt
     23 mekanism
     12 mekanismen
     45 mekanismer
     12 mekanismerna
      1 mekanistiska
      1 mekonium
      2 mekoniumet
      1 mekoniumfärgat
      1 mel
     17 melamin
      2 melaminet
      3 melaminplast
      2 melaminskandalen
      1 melampos
      1 melancholie
      1 melanesians
      1 melanesiskt
      3 melanie
     10 melanin
      2 melaniner
      1 melaninfläckar
      1 melanininnehållande
      1 melaninkoncentrerande
      1 melanism
     31 melankoli
      2 melankolier
      4 melankoliker
      7 melankolikern
      1 melankolikerns
      4 melankolin
      3 melankolisk
      5 melankoliska
      1 melanocortinreceptor
      3 melanocyter
      2 melanocyterna
      2 melanom
      1 melasma
     33 melatonin
      1 melatoninproduktionen
      1 melbourne
      1 melbournes
      1 melena
      1 melia
      1 melinda
   1055 mellan
      2 mellanamerika
      1 mellanavstånd
      1 mellanbarn
      1 mellanblödningar
      1 mellandos
      1 mellaneuropa
      1 mellaneuropeiska
      1 mellanfas
      1 mellanformer
      2 mellanfotsben
      1 mellangården
      1 mellangärdesnerven
      5 mellangärdet
      1 mellanhänder
      9 mellanhjärnan
      1 mellanhjärnans
      1 mellanlager
      1 mellanlägg
      4 mellanliggande
      2 mellanmänskliga
      1 mellanolja
      5 mellanörat
      1 mellanöreinflammation
      1 mellanöron
     10 mellanöstern
      1 mellanprodukt
      1 mellanregistret
     19 mellanrum
      1 mellanrummet
      2 mellanrumsborstar
      6 mellanrumsborste
      1 mellanrumsborsten
      1 mellanskikt
      1 mellanskiktet
      1 mellanstation
      1 mellanstatliga
      5 mellansteg
      2 mellanstegen
      1 mellanstora
      1 mellanstycke
      1 mellanstycket
      1 mellansubstans
      1 mellansvår
      2 mellansverige
      3 mellanting
      1 mellanvåg
      2 mellanväggen
      5 mellanvärd
      1 mellanvärdar
      1 mellea
     12 mellersta
      8 mellitus
      1 melodin
      1 melodislinga
      1 melos
      1 melville
      1 melvilleöarna
      2 memantin
      1 member
     26 membran
      2 membranbundna
      1 membrandelar
      2 membrandelen
      1 membraner
     10 membranet
      1 membranets
      1 membranfilter
      1 membrankanaler
      1 membranomsluten
      1 membranomslutna
      2 membranpotential
      5 membranpotentialen
      2 membranprotein
      1 membranstörande
      3 memento
      1 memorerar
      2 memorial
      1 memory
   2447 men
      4 mena
     26 menade
      1 menades
      1 menafrivac
     95 menar
     12 menarche
      1 menarchen
     29 menas
      7 menat
      2 mendel
      1 mendelejevs
      1 mendor
      1 menevis
      1 mengele
      1 meng�mok
      1 menigheten
      1 menigokocksjukdom
     35 mening
     11 meningar
      1 meningeal
      2 meningeala
     14 meningen
      8 meningeom
      1 meningierna
      3 meningiom
      1 meningioma
      1 méningiome
    118 meningit
      3 meningitbältet
      6 meningiten
      1 meningitfall
      1 meningitidesgrupperna
      4 meningitidis
      1 meningitidishaemophilus
      1 meningitis
      3 meningocele
      1 meningococcus
      2 meningokock
      1 meningokockepidemier
     10 meningokocker
      1 meningokockgrupp
     10 meningokockmeningit
      4 meningokocksjukdom
      1 meningokockvacciner
      2 meningovaskulär
      4 meningsfull
      2 meningsfulla
      7 meningsfullhet
      1 meningsfullheten
      7 meningsfullt
      2 meningslös
      3 meningslöst
      1 meningsmotståndare
      1 meningsskapande
      1 menisk
      2 menkes
      1 menlig
      1 mennarke
      1 mennesket
      1 menninger
      1 menningerkliniken
      9 menopaus
      8 menopausen
      1 menorragi
     15 mens
      3 mensa
      1 mensbesvär
      2 mensblod
      2 mensblodet
      1 mensblödning
      5 menscykel
      8 menscykeln
      1 mensdebut
      3 mensen
      1 mensens
      2 mensis
     10 menskopp
     10 menskoppar
      1 menskopparna
      9 menskoppen
      1 menskoppsanvändning
     16 mensskydd
      1 mensskyddet
      1 menstruaionscykeln
      1 menstruaitonspsykos
      1 menstrualis
     29 menstruation
     29 menstruationen
      3 menstruationens
      4 menstruationer
      4 menstruationerna
      3 menstruationsblod
      5 menstruationsblodet
      2 menstruationsblödningar
      2 menstruationsblödningen
      7 menstruationscykel
     25 menstruationscykeln
      1 menstruationsdebut
      2 menstruationsliknande
      1 menstruationsmönstret
      1 menstruationsperioden
      5 menstruationspsykos
      6 menstruationspsykoser
      1 menstruationsrubbningar
      1 menstruationsskydd
      1 menstruationssmärta
     11 menstruationsstörningar
      1 menstruationsvätska
      1 menstruerande
      1 menstruerar
      4 mensvärk
      1 mensvärken
      1 mensvärksliknande
      1 mentagrophytes
     54 mental
     31 mentala
      1 mentalhälsolagstiftning
      1 mentalhälsolagstiftningen
      1 mentalhygien
      1 mentalisera
      1 mentaliseringsförmåga
      1 mentalsjukdom
      3 mentalsjukdomar
      1 mentalsjukdomarna
      3 mentalsjukhus
      3 mentalsjukhusen
      1 mentalsjukhuset
      1 mentalsocial
     12 mentalt
      2 mentalvården
      1 mentalvårdslagstiftning
      3 mentol
      2 mentor
      1 mentorer
      1 mentorn
    897 mer
    133 mera
      1 merci
      2 merck
      1 mercoire
      1 mercurialis
      1 mercurius
      2 mercury
      1 mercyful
      1 merely
      1 merendera
      1 merengue
      1 meridianer
      1 meridianpunkter
      2 mering
      1 merings
      1 meripilus
      1 merkantilismen
      1 merkaptaner
      1 merkostnadslån
      1 merle
      1 merlegen
      1 merlin
      1 meroencefali
      1 meropenem
      2 merozoiter
      1 merozoiterna
      7 merparten
      2 merricks
      1 merrit
      5 mesalazin
      1 mesangialceller
      1 mescal
      1 mescalråvara
      1 mesencephalon
      1 mesenchymala
      1 mesenkymala
      1 mesenkymatisk
      1 mesenterium
      5 mesh
      2 meshtermer
      1 meskalin
      3 mesmer
      1 mesna
      1 mesocefal
      1 mesoderm
      1 mesodermet
      2 mesogloea
      1 mesokortikala
      2 mesolimbiska
      2 mesopotamien
      1 mesotel
      5 mesoteliom
      5 mesotheliom
      1 mesotheliomets
      1 messias
      2 messina
    273 mest
     33 mesta
      8 mestadels
      1 metaamfetamin
      4 metaanalys
      1 metaanalysartikel
      7 metabol
     13 metabola
      2 metaboliserar
      4 metaboliseras
      1 metaboliserat
      3 metabolisk
     14 metaboliska
     23 metabolism
      5 metabolismen
      1 metabolistiska
      2 metabolit
      1 metaboliten
      9 metaboliter
      3 metaboliterna
     10 metabolt
      1 metaborater
      3 metaborsyra
      1 metabotropa
      1 metadioxidifenylamin
      2 metadon
      1 metadonbussar
      3 metafor
      1 metaforen
      1 metafysik
      1 metafysiken
      5 metafysisk
      1 metafysiska
     30 metall
      2 metallbågar
      1 metallbygel
      1 metallclips
      1 metalldelar
      1 metallegering
      1 metallegeringar
      5 metallen
      1 metallens
     12 metaller
      2 metallerna
      1 metallernas
      1 metallers
      1 metallföreningar
      1 metallgjuterier
      2 metallisk
      1 metalliska
     12 metalliskt
      1 metallkant
      1 metallkärl
      1 metallkatalysator
      1 metallklämma
      3 metallnät
      1 metalloproteinaser
      1 metallotionein
      1 metallplattor
      1 metallring
      2 metallrör
      1 metallsalter
      1 metallsalterna
      1 metallsmak
      1 metallspadar
      1 metallspeglar
      1 metallstag
      1 metallstycke
      1 metallstycken
      4 metalltråd
      1 metalltrådar
      1 metalltråden
      1 metalltuben
      1 metallurgiska
      1 metallurgiskt
      1 metallvärde
      1 metallvärdet
      1 metallvaror
      1 metallverk
      1 metallverktyg
      1 metallyta
      1 metallytad
      1 metallytan
      5 metamfetamin
      2 metamina
      1 metamorf
      1 metamorfa
      1 metamorfism
      1 metamorfismprodukt
      5 metamorfos
      1 metamyelocyten
      5 metan
      1 metanal
      1 metangas
      1 metangasframställning
     21 metanol
      1 metanolförgiftning
      1 metansyra
      4 metaplasi
      2 metaplasier
      2 metapneumovirus
      1 metastabila
      5 metastas
     27 metastaser
      5 metastasera
      2 metastaserad
      3 metastaserande
      6 metastaserar
      1 metastaseras
      1 metastaserat
      1 metastaserats
      3 metastasering
      1 metastaseringsplatser
      3 metastaserna
      1 metastatiska
      7 metastudie
      3 metastudier
      1 metateorin
      2 metenamin
      3 meteorism
     78 meter
      1 meterhög
      1 meterhöga
      1 meterlång
     10 meters
      1 metervara
      3 metformin
      2 methemoglobin
      1 methemoglobinemi
      2 method
      1 methods
      2 methusalem
      1 methylhexenoic
      2 meticillin
      2 meticillinresistens
      1 meticillinresistent
      4 meticillinresistenta
      1 métiers
    168 metod
    143 metoden
      3 metodens
    173 metoder
      1 metoderhjälpmedel
     21 metoderna
      1 metodernas
      3 metodik
      2 metodiken
      1 metodiska
      1 metodiskt
      4 metodologiska
      1 metodstyrd
      5 metotrexat
      1 metoxykatekolaminer
      4 metrik
      1 metron
      5 metronidazol
      1 metropolitan
      1 metyl
      1 metylalkohol
      2 metylamfetamin
      1 metylbromid
      1 metylcyanoakrylat
      1 metylcyanopropenoat
      3 metyldopa
      1 metylenblått
      1 metylendiresorcin
      1 metylenklorfluorid
      1 metylepoxioktadekan
      1 metylergometrin
      1 metylergometrintartrat
      1 metylering
      3 metylfenidat
      1 metylfenol
      1 metylgrupp
      1 metylimidazol
      1 metylisopropylfenol
      1 metyljodid
      1 metylketoner
      1 metylklordifluorid
      1 metylklorid
      1 metylkvicksilver
      1 metylmetkatinon
      1 metylparaben
      1 metylpropanol
      1 metylsalicylat
      1 metyltetrametyltrimetylsilyloxydisiloxanylpropyl
      1 metylumbelliferon
      2 mev
      1 mexicanum
      6 mexico
      2 mexikansk
      1 mexikanska
      1 mexikanskt
     15 mexiko
      2 meyer
      4 meyers
      1 meyersmits
      1 mezerein
      1 mezereum
      1 mezeriyn
      1 mezerum
      1 mezger
      1 mfd
     13 mfl
      1 mfp
     37 mg
      1 mgdag
      2 mgdl
      1 mgfealalsioohho
      1 mgkg
      2 mgl
      3 mgml
      1 mgohsio
      1 mgvecka
      1 m�h
      1 mha
      6 mhc
      1 mhcalleler
      2 mhckomplex
      1 mhckomplexen
      1 mhcmolekyler
      1 mhcstrukturer
      1 mhydrokinon
      2 mhz
      1 miasajter
      1 miasm
      3 miasmer
      1 miasmhypotes
      1 miasmteori
      1 miasmteorin
      1 mic
      1 micellkoncentration
     16 michael
      1 michail
      1 michaut
      2 michel
      1 michelangelo
      1 michele
      1 michelle
      1 michigan
      1 michio
      1 microarrays
      1 microcefali
      1 microcephala
      1 microcid
      1 microflora
      1 microlax
      1 microlepidotus
      1 microneurokirurgin
      1 microplus
      1 microsporum
      1 microti
      1 microtubilii
      1 microtubuli
      1 midaxillarlinjen
      2 midazolam
      2 middagar
      1 middagsgästerna
      1 middagshöjd
      1 middagstiden
      1 middle
      1 mideighteenthcentury
      7 midja
      6 midjahöftkvot
      2 midjahöftkvoten
     10 midjan
      1 midjans
      1 midjebälte
      8 midjemått
      3 midjemåttet
      1 midjeomfång
      1 midjeväska
      1 midnfulnessbaserad
      1 midsommar
      1 midsommarblomster
      1 midsommardagen
      1 midsommartid
      2 miele
      9 mig
     18 migrän
      4 migrans
      1 migrating
      1 migration
      1 migrera
      2 migrerande
      2 migrerar
      1 migrerat
      1 mike
      2 mikro
      1 mikroadenom
      2 mikroakupunktur
      1 mikroampere
      1 mikroangiopati
      1 mikrob
      1 mikroba
      8 mikrober
      2 mikroberna
      1 mikrobiell
      2 mikrobiella
      1 mikrobiologen
      6 mikrobiologi
      1 mikrobiologins
      2 mikrobiologisk
      3 mikrobiologiska
      1 mikrobiska
      5 mikrocefali
      1 mikrocytär
      1 mikrofloran
      6 mikrofon
      1 mikrofonen
      1 mikrofoner
      8 mikroftalmi
      1 mikrogamofyten
      1 mikrogliaceller
      6 mikrogram
      1 mikrograml
      1 mikroinplantat
      1 mikrokeratom
      1 mikrokirurgi
      1 mikrokocker
      1 mikrokolonier
      1 mikrokosmos
      1 mikrokretsar
      1 mikrolavemang
      1 mikromatrisanalys
      1 mikromatrisanalyser
      2 mikromatriser
      1 mikrometastaser
     12 mikrometer
      1 mikromiljö
      2 mikromiljön
      1 mikromoll
      2 mikronäringsämnen
      5 mikroorganism
      2 mikroorganismen
     69 mikroorganismer
      8 mikroorganismerna
      3 mikroorganismernas
      1 mikroorganismers
      1 mikropartiklar
      2 mikropenis
      1 mikropyle
      1 mikrosimulering
     24 mikroskop
      1 mikroskopet
      3 mikroskopi
      6 mikroskopisk
     15 mikroskopiska
      2 mikroskopiskt
      1 mikroskopundersökning
      1 mikrosomala
      2 mikrosvampar
      1 mikrosvampars
      1 mikrosystem
      1 mikrotabletter
      1 mikrotabletterna
      1 mikrotom
      1 mikrotromboser
      1 mikrotubuli
      3 mikrovågor
      6 mikrovågsugn
      1 mikrovaskulär
      1 mikrovaskulära
      5 mikrovilli
      1 mikrovilliutskott
      1 miktera
      2 miktion
      1 miktionsfrekvens
      1 miktionsuretrocystografi
      2 mil
      1 milan
     24 mild
      9 milda
     18 mildare
      2 mildra
      1 mildrabota
      1 mildrar
      5 miliaria
      4 miliartuberkulos
      1 milier
      6 militär
     14 militära
      1 militärbaracker
      1 militärbårar
      1 militärbasen
      2 militären
      1 militärens
      2 militärer
      1 militärflygplan
      1 militärläkare
      1 militärpolis
      5 militärt
      2 militärtjänst
      4 miljard
      1 miljardbelopp
      1 miljarddel
     26 miljarder
      1 miljarderusd
     76 miljö
      1 miljöaktivister
      1 miljöändringar
      1 miljöarbete
      2 miljöaspekter
      1 miljöåtgärder
      2 miljöbalken
      2 miljöbrott
      1 miljöchef
      3 miljöeffekter
     35 miljöer
      1 miljöerna
      1 miljöfaktor
     17 miljöfaktorer
      3 miljöfaktorers
      1 miljöfarlig
      5 miljöfarliga
      1 miljöfarlighetsbedömning
      1 miljöfarlighetssymbol
      1 miljöfarligt
      2 miljöförändringar
      1 miljöförstöring
      1 miljöförstöringen
      4 miljögift
      8 miljögifter
      1 miljögiftet
      1 miljöinformation
      1 miljöinsatser
      1 miljöklassad
      1 miljömärkningarna
      1 miljömässig
      6 miljömässiga
      1 miljömässigt
      5 miljömedicin
      1 miljömedicinsk
      1 miljömedicinska
     18 miljon
     51 miljön
      1 miljönämnden
    158 miljoner
      2 miljöns
      5 miljontals
      1 miljöorsakad
      1 miljööverdomstolen
      1 miljöpartiet
      2 miljöpåverkan
      5 miljöproblem
      1 miljöprogram
      1 miljörelaterade
      1 miljörisker
      1 miljörörelsen
      1 miljörörelser
      1 miljösamordnare
      1 miljöskadligt
      2 miljöskador
      1 miljöskadorna
      4 miljöskäl
      1 miljösynpunkt
      1 miljöutskott
      1 miljöval
      1 miljövänliga
      1 miljövänligare
      3 miljövänligt
      1 miljövård
      1 milkshake
      1 millenniedeklarationen
      1 millenniemål
      4 millenniemålen
      1 millennieskiftet
      1 millennietoppmötet
      2 miller
      1 millerblad
      1 milleri
      8 milligram
      8 milliliter
     31 millimeter
      1 millimeterbreda
      1 millimeters
      1 millimetertjocka
      1 millisievert
      1 millivolt
      1 mills
      1 milstolpar
      1 milstolpe
     10 milt
      2 milton
      1 milwaukee
      1 milwaukeeprotokollet
      1 mimicry
      1 mimik
      1 mimiken
      1 mimos
      8 min
      1 mina
      2 mind
      1 minderåriga
      1 mindervärda
      3 mindfulness
      3 mindfulnessbaserad
    505 mindre
      1 minelli
     18 mineral
      1 mineralämnen
      1 mineralbrist
      1 mineralbrister
     17 mineraler
      1 mineralerna
      5 mineralet
      1 mineralfiber
      1 mineralförening
      1 mineralförgiftning
      2 mineralglas
      1 mineralgrupperna
      1 mineralkortikoidreceptorer
      1 mineralnamnet
      1 mineralog
      1 mineralogi
      1 mineralolja
      1 mineralpreparat
      1 mineralriket
      2 mineralsalter
      2 mingdynastin
      1 mini
      1 miniatyr
      1 miniatyrisering
      1 minibussar
      1 minifom
      1 minikamera
      1 minikurs
      7 minimal
      2 minimala
      2 minimalinvasiva
      2 minimalt
     16 minimera
      4 minimerar
      2 minimeras
      1 minimienergin
      1 minimikraven
      1 minimizer
      1 minimizerbh
      4 minimum
      1 minimumintensity
      5 minipiller
      1 minister
      1 ministerium
      1 ministrar
      1 minitampong
      1 minitrauma
      2 mink
      1 minkfarmar
      1 minkowski
      1 minkowskis
      1 minmera
      1 minnas
     26 minne
     13 minnen
      1 minnesbilder
      1 minnesbildning
      1 minnesceller
      1 minnesfel
      5 minnesförlust
      1 minnesförluster
      1 minnesförmåga
      1 minnesformering
      1 minnesfunktion
      1 minnesfunktionen
      1 minnesfunktioner
      1 minnesgåva
      1 minneskapaciteten
      1 minneslek
      1 minneslucka
      2 minnesmetall
      1 minnesmetallen
      1 minnesmetaller
      1 minnesoscilloskop
      1 minnesota
      1 minnesotamodellen
      1 minnesplast
      1 minnesprestationer
      5 minnesproblem
      1 minnesprocessen
      1 minnesskärm
      5 minnesstörningar
      3 minnessvårigheter
     13 minnet
      8 minns
      1 minoiska
      3 minor
      1 minora
     11 minoritet
      2 minoriteten
      2 minoriteter
      1 minoriteterna
      1 minoritetsgrupperna
      1 minoritetssamhällen
    217 minska
     83 minskad
     35 minskade
      2 minskades
      3 minskande
    174 minskar
     24 minskas
     47 minskat
      1 minskaundvika
     21 minskning
      8 minskningen
      1 minspel
    152 minst
     32 minsta
      1 minstbakterier
      2 mint
      5 minus
      1 minusgrader
      1 minuspol
      1 minussträngad
      1 minusvärden
     36 minut
      3 minute
      2 minuten
     64 minuter
      1 minuterna
      5 minuters
      1 minutertimmar
      2 minutvolym
      3 minutvolymen
      2 mios
      1 miosis
      2 mip
      2 mirabilia
      1 miracidier
      2 mirakelkurer
      1 mirakelmedicin
      1 mirakelmedicinen
      1 mirakelmediciner
      1 mirakelpiller
      1 mirakulösa
      1 mircea
      2 mirescu
      1 mirror
      3 misär
      1 miskar
      2 mismeasure
      1 miso
      1 mison
      2 misophonia
      4 misosoppa
      2 misosoppan
      4 miss
      1 missa
      1 missade
      1 missar
      1 missas
      1 missat
      1 missbedömd
      1 missbelåtenhet
      4 missbildade
     30 missbildning
     36 missbildningar
      1 missbildningarna
     10 missbildningen
      1 missbildningens
      2 missbildningsbenäget
      1 missbildningssyndrom
      1 missbildningstumör
     53 missbruk
      1 missbruka
      3 missbrukar
     13 missbrukare
      2 missbrukaren
      1 missbrukarledet
      1 missbrukarnas
      5 missbruket
      1 missbrukets
      2 missbruks
      1 missbrukskarriär
      1 missbrukskategorier
      1 missbruksmedel
      1 missbruksproblem
      1 missbrukspsykiatri
      1 missbruksrisk
      1 missbruksrisken
      1 missbrukssyfte
      2 missbruksutredningen
      2 missbruksvård
      1 missbruksvården
      2 missed
     44 missfall
      3 missfallet
      2 missfärga
      1 missfärgad
      1 missfärgade
      1 missfärgande
      1 missfärgas
      1 missfärgat
      7 missfärgning
      2 missfärgningar
      2 missfärgningen
      1 missformat
      1 missformningar
      4 missförstånd
      1 missförstått
      1 missförståtts
      2 missfoster
      1 missgärningsbalken
      1 missgestaltande
      1 missgynna
      1 missgynnad
      1 missgynnas
      2 misshagliga
      6 misshandel
      1 missiler
      1 missionären
      1 mississippideltat
      1 mississippinew
      1 misskötande
      1 missleda
      1 missledande
      4 misslyckad
      2 misslyckade
      1 misslyckades
      6 misslyckande
      3 misslyckanden
      8 misslyckas
      1 misslyckat
      7 misslyckats
      1 missnöjd
      1 missnöjdhet
      1 missnöje
      1 missnöjet
      1 missöden
      1 missos
      2 missouri
     10 misstag
      1 misstänka
      4 misstankar
      1 misstankarna
      7 misstänkas
     25 misstanke
      1 misstanken
      7 misstänker
     17 misstänks
      8 misstänksamhet
      1 misstänksamma
      1 misstänksamt
     22 misstänkt
     14 misstänkta
      2 misstänkte
      2 misstänktes
      6 misstas
      2 misstolka
      1 misstolkar
      1 misstolkas
      1 misstolkningar
      1 misstror
      1 misstycker
      1 missummarsurta
      2 missuppfattas
      5 missuppfattning
      1 missuppfattningen
      1 missväxt
     18 missvisande
      4 miste
      1 mister
      1 mitchells
      3 mitella
      3 mithridat
      7 mithridates
      1 mithridatet
      1 mithridatets
      1 mithridatica
      1 mithridaticum
      1 mitogen
      1 mitokondriella
      1 mitokondriellt
      9 mitokondrier
      3 mitokondrierna
      1 mitokondriernas
      1 mitokondriskt
      5 mitos
      1 mitoser
      1 mitotiska
      1 mitralis
      3 mitralisklaffen
      1 mitridat
     21 mitt
      2 mittemellan
     65 mitten
      1 mittentån
      1 mittersta
      9 mitthjärnan
      3 mittlinjen
      2 mittnerv
      1 mittpartibr
      1 mittportionsprov
      1 mittpunkt
      1 mitträcke
      1 mittremsa
      2 mittremsan
      1 mittstjälken
      1 mittsträng
      1 miva
      1 mixers
      2 mixtur
      1 mixturen
      1 mj
      9 mjäll
      1 mjällbildning
      1 mjällproduktionen
     14 mjältbrand
      1 mjältbrandsattackerna
      1 mjältbrandsbakterier
      1 mjältbrandsbakterierna
      1 mjältbrandsutbrott
     11 mjälte
     16 mjälten
      6 mjöl
      4 mjöldagg
      1 mjöldaggssvamparna
      1 mjöldaggssvampen
     20 mjöldryga
      2 mjöldrygan
      1 mjöldrygeepidemi
      4 mjöldrygeförgiftning
      1 mjöldrygeförgiftningar
      1 mjöldrygeinfekterad
      1 mjöldrygeinfektion
      2 mjöldrygesvampen
      1 mjöldrygorna
      2 mjölet
      1 mjölig
     53 mjölk
      1 mjölkade
      1 mjölkaktigt
      4 mjölkallergi
      1 mjölkallergiker
      1 mjölkallergiska
      2 mjölkavsöndringen
      1 mjölkbaserad
      1 mjölkbildande
      1 mjölkbildning
      1 mjölkcisternen
      1 mjölkdrickande
     12 mjölken
      2 mjölkersättning
      1 mjölkersättningar
      1 mjölkerskor
      1 mjölkfettet
      1 mjölkflödet
      1 mjölkgång
      1 mjölkgångar
      5 mjölkgångarna
      1 mjölkgångsepitel
      1 mjölkgångsröntgen
      1 mjölkhaltig
      1 mjölkiga
      2 mjölkkanalerna
      1 mjölkkartong
      1 mjölkkobesättningar
      2 mjölkkor
      1 mjölkkörtel
      1 mjölkkörtlar
      5 mjölkkörtlarna
      1 mjölkkörtlarnas
      2 mjölkmaskiner
      3 mjölkning
      1 mjölkningspersonalen
      1 mjölkorganet
      1 mjölkpigor
      1 mjölkproducerande
     13 mjölkprodukter
      1 mjölkprodukters
      3 mjölkproduktion
      2 mjölkproduktionen
      1 mjölkprotein
      1 mjölkproteiner
      1 mjölkpulver
      2 mjölksaft
      2 mjölksaften
      1 mjölksekretion
      5 mjölkskorv
      1 mjölkskorven
      4 mjölksocker
      7 mjölkstockning
      2 mjölkstockningen
      1 mjölkstockningens
      9 mjölksyra
      1 mjölksyrabakterier
      1 mjölksyrabakterierna
      1 mjölksyran
      1 mjölksyratröskeln
      1 mjölksyrebakterier
      1 mjölksyror
      1 mjölktänder
      1 mjölkutsöndring
      1 mjölliknande
      1 mjölproducerande
      1 mjölskivling
      1 mjölskivlingen
      1 mjölsorter
      1 mjuddelsabscesser
     20 mjuk
     29 mjuka
      3 mjukar
      6 mjukare
      3 mjukas
      6 mjukdelar
      1 mjukdelarna
      1 mjukdels
      2 mjukdelsinfektioner
      1 mjukglass
      2 mjukgöra
      6 mjukgörande
      3 mjukgörare
      1 mjukhet
      1 mjukmedel
      1 mjukna
      1 mjuknar
      1 mjuknat
      1 mjukost
      3 mjukpapper
      1 mjukpappersprodukterna
      2 mjukplast
      1 mjukröntgenstrålning
     10 mjukt
      3 mjukvara
      1 mjukvaran
      1 mjukvaruföretag
      2 mjukvävnad
      1 mjukvävnader
      6 mkomponent
      3 mkomponenten
      1 mkomponenter
      1 mkopp
      1 mkubikmeter
     30 ml
      1 mldygn
      1 mlkgh
      2 mlkgmin
      1 mlkg�min
      1 mlmin
     97 mm
      2 �mm
      2 mma
      4 mmc
      1 mmcd
      1 mmhg
      2 mmode
      7 mmoll
      2 mmp
      1 mmt
      4 mno
      1 mnsblodgruppssystemet
      1 mnssystemet
      4 mo�ambique
      1 mobbare
      4 mobbing
      3 mobbning
      1 möbel
      1 möbelmässan
      1 möbeltassar
      1 mobil
      2 mobila
      1 mobilen
      1 mobilfas
      4 mobilisera
      2 mobiliserande
      4 mobilisering
      1 mobiliseringen
      1 mobilitas
      1 mobility
      1 mobilkamera
      1 mobillyftar
      7 mobiltelefon
      1 mobiltelefonanvändning
      5 mobiltelefoner
      1 mobiltelefoners
      1 mobiltelefonföretag
      1 mobiltelefonsignaleroch
      4 möbler
      1 moby
      2 mockasinsvamp
      1 mod
      2 modafinil
      4 modaliteter
      1 mödan
     12 mode
      1 modedesignern
      3 modehusen
      1 modeindustrin
      1 model
     19 modell
      9 modellen
      1 modellens
     22 modeller
      1 modelleras
      2 modellering
      7 modellerna
      3 modellinlärning
      1 modellr
      1 modemedvetna
      1 modeplagg
      7 moder
      4 moderat
      2 moderator
      1 moderatormaterial
      1 moderbolag
      1 moderbolagets
      2 modercell
      1 moderindividen
      1 moderinstinkter
      1 moderkaka
     18 moderkakan
      2 moderkakans
      2 moderkorset
      1 moderlivet
    113 modern
     99 moderna
      8 modernare
      1 modernhan
      1 moderniseringar
      1 moderniseringen
      3 modernitet
     16 moderns
      7 modernt
      1 moderorganisation
      1 moderplantan
      1 moderrelationen
      1 moderrullarna
      1 moders
      3 modersbeteenden
      1 moderskänslor
      1 moderskänslorna
      3 modersmål
      4 modersmjölk
      2 modersmjölken
      1 modersmjölkersättning
      1 modersmjölksersättningar
      1 modersubstans
      1 modersvulsten
      1 modertumören
      1 modeskaparna
      1 modesta
     12 modet
      2 modetillbehör
      1 modification
      5 modifiera
      1 modifierad
      9 modifierade
      1 modifierades
      1 modifierande
      3 modifierar
      5 modifieras
      3 modifierat
      2 modifiering
      1 �modifikation
      3 modifikationer
      1 modifying
      2 mödomshinnan
      1 mödosamt
      2 mödradödlighet
      3 mödrahälsovård
      1 mödrahälsovården
     28 mödrar
      2 mödrarna
      2 mödrarnas
      1 mödrars
      3 mödravård
      5 mödravården
      2 mödravårdscentral
      1 mödravårdsmottagningen
      1 mods
      3 moduco
      2 modul
      1 modulärt
      1 modulationsteorin
      1 modulera
      2 modulerar
      1 modulerare
      3 moduleras
      2 moduleringar
      1 mody
      8 mögel
      1 mögelbildningen
      1 mögelsläktet
      2 mögelsporer
      1 mögelsvamp
      7 mogen
      5 moget
      1 möglet
      1 möglets
      1 möglig
      1 mögliga
      1 mögligt
     22 mogna
      5 mognad
      3 mognaden
      1 mognadsfråga
      2 mognadsgrad
      1 mognadsprocess
      1 mognadsprocessen
     15 mognar
      2 mognat
      1 mogulriket
      2 moh
      1 mohs
      1 mojito
     34 möjlig
     45 möjliga
      1 möjligaste
     42 möjligen
      2 möjliggjorde
      1 möjliggjordes
      1 möjliggjort
      2 möjliggjorts
     17 möjliggör
     11 möjliggöra
      3 möjliggörs
     76 möjlighet
     33 möjligheten
     25 möjligheter
      9 möjligheterna
    177 möjligt
      3 möjligtvis
      1 mök
      1 mokasen
      2 moksha
      3 mola
      2 molagraviditet
      1 molarerna
      1 molekulära
      1 molekyer
     23 molekyl
      8 molekylär
      6 molekylära
      2 molekylärbiologi
      1 molekylärbiologin
      1 molekylärbiologins
      1 molekylärbiologisk
      2 molekylärbiologiska
      1 molekylärdiagnostik
      1 molekylärt
     14 molekylen
      1 molekylens
     48 molekyler
      9 molekylerna
      1 molekylernas
      2 molekylers
      1 molekylformeln
      1 molekylmassan
      1 molekylsönderdelande
      1 molekylvikt
      1 molekylvikten
      3 moleler
      1 molift
      1 moli�re
      3 moll
      1 mollaretmeningit
      1 mölle
      1 mollusker
      2 molmassa
      2 moln
      1 mölnlycke
      1 molnsådd
      1 molotovcocktails
      1 molvolym
      3 molybden
      1 molybdenmalm
      6 moment
      3 momentant
      1 momentet
      1 moms
      1 momsbefriat
      1 momsplitktigt
      1 monaminerga
      1 mondeville
      1 monel
      1 mongoler
      3 mongolerna
      1 mongolfläck
      3 mongolfläcken
      1 mongolism
      1 mongoloid
      1 monica
      1 monika
      1 monila
      1 monilia
      1 moniliformis
      1 monitor
      2 monitoring
      2 moniz
      1 monkliniska
      1 monoaddukt
      2 monoaddukter
      1 monoaminer
      1 monoaminoxidas
      1 monobaktamer
      1 monobutyltenn
      2 monocytär
      1 monocytära
      3 monocyter
      1 monocytogenes
      1 monoetylenglykol
      1 monofluoridfosfat
      3 monogama
      1 monogen
      1 monogenea
      1 monografi
      1 monografier
      1 monografin
      2 monogram
      1 monohydratet
      1 monohydratets
      1 monoik
      1 monojodtyrosin
      1 monokarp
      2 monokarper
      2 monokel
      2 monokeln
      2 monokini
      1 monokinin
      1 monoklar
      3 monoklint
      2 monoklonal
      7 monoklonala
      1 monoklonalt
      1 monokromatisk
      1 monolog
      2 mononegavirales
      1 mononeuropatier
      1 mononukleära
      2 mononukleos
      3 monopol
      1 monorkism
      1 monos
      1 monosackarid
      2 monosackariden
      3 monosackarider
      1 monosodiumglutamat
      1 monosomi
      1 monosomier
      1 monosubstituerade
      1 monosynaptisk
      2 monoteistiska
      3 monoterapi
      1 monoton
      3 monotona
      1 monotont
      2 monotypiska
      2 monsanto
      1 monsantoprocessen
      5 monster
     28 mönster
      1 mönsterbildande
      1 mönsterigenkänning
      1 mönsterstickades
      1 mönstertryck
      1 mönstra
      2 mönstrad
      1 mönstrade
      2 mönstrat
      2 monstret
      4 mönstret
      1 monstrosus
      1 montagearbete
      3 montagnier
      1 montagniers
      1 montagu
      2 montaguadalen
      2 montana
      1 montelukast
      1 montenier
      1 monterad
      4 monterade
      1 monterar
      6 monteras
      1 monterats
      3 montering
      1 monteringar
      1 montezumas
      1 montgomerys
      1 montignac
      2 montignacdieten
      1 montmartre
      1 montparnasse
      1 montpellier
      3 montrealprotokollet
      1 monumentala
      1 moon
      3 moped
      1 mopedförare
      3 mopedister
     17 mor
      1 mora
      1 moraknivskirurgi
      8 moral
      4 moralisk
      5 moraliska
      1 moralisketisk
      4 moraliskt
      2 moralism
      1 moralistiska
      1 morallagar
      2 moraxella
      1 morbarn
      2 morbiditet
      2 morbilli
      2 morbillisläktet
      1 morbillivirus
      1 morborum
      3 morbus
      1 mörby
      5 mord
      1 mördade
      1 mördar
      1 mördarceller
      3 mördare
      2 mördat
      1 mordbrand
      1 mordet
      2 mordoffer
      1 mordraseri
      1 mordutredning
      1 morement
      1 morfar
      3 morfem
      1 morfematisk
      1 morfematiskt
      1 morfematisktskt
      1 morfemgränser
     11 morfin
      1 morfinbruk
      1 morfinet
      1 morfininjektioner
      1 morfinism
      8 morfologi
      1 morfologin
      1 morfologiska
      3 morfologiskt
      1 morgagni
      1 morgan
      1 morgnar
      1 morgnarna
      9 morgon
     19 morgonen
      1 morgonstånd
      1 morgonstela
      1 morgontemperatur
      1 morgontrötthet
      1 mori
      1 morihei
      1 moriska
      1 moritz
     10 mörk
     11 mörka
     29 mörkare
      1 mörkblå
      3 mörkbrun
      2 mörkbrunt
      6 mörker
      1 mörkerseende
      1 mörkerseendet
      2 mörkertal
      4 mörkertalet
      1 mörkfältsmikroskopi
      1 mörkfärgning
      2 mörkfjälliga
      1 mörkgrön
      1 mörkgröna
      1 mörkgula
      1 mörkhåriga
      2 mörkhyad
      2 mörkhyade
      1 mörklagts
      1 mörklila
      1 mörkna
      1 mörknar
      1 mörkret
      1 mörkröda
     12 mörkt
      1 mormorsglasögonen
      1 mormorsmor
      1 mörner
      1 morötter
      1 morphy
      1 morrison
      1 mörsil
      1 morsuvae
     13 mortalitet
      9 mortaliteten
      1 mortelstötar
      1 mortem
      1 morten
      2 morton
      2 mortons
      1 morula
      2 morulan
      1 mos
      1 mosaicism
      1 mosaicistisk
      1 mosaicistiska
      1 mosaikism
      2 mosaiska
      1 mosby
      1 moseböcker
      2 mosebok
      5 moseboken
      1 mosebokens
      1 moseleys
      1 moseleyum
      1 moshe
      2 moskitfisk
      3 moskva
      1 mosley
      2 mosonmagyaróvár
     30 möss
      1 mossa
      1 mössa
      1 mossar
      1 mösseberg
      3 mössmärke
      2 mossor
      1 mössor
      1 most
   1286 mot
     10 möta
      1 motalahäxan
      4 mötande
      2 motang
      1 motangrepp
      1 motantibiotika
      2 motarbeta
      1 motarbetade
      2 motarbetas
      1 motåtgärd
      1 motåtgärder
      2 motbevisa
      7 motbevisad
      2 motbjudande
      7 möte
      9 möten
      4 mötena
      7 möter
      1 moterneuronskador
      1 mötes
      7 mötet
      3 motgångar
      7 motgift
      1 motgiftet
      2 mothäxor
      1 mother
      2 motila
      2 motilitet
      1 motilitetsgrad
      1 motilitetsgraden
     29 motion
      2 motioner
      4 motionera
      1 motionmedierad
      1 motionsförbud
      1 motionslokaler
      1 motionsträning
      2 motionsvanor
      9 motiv
     14 motivation
      4 motivationen
      1 motivationssystem
      1 motivbilderna
      5 motiven
      4 motivera
      4 motiverad
      3 motiverade
      2 motiverades
      2 motiverande
      3 motiverar
      7 motiveras
      3 motivering
      2 motiveringen
      1 motivet
      1 motjoner
      1 mötley
      3 motmedel
     10 motor
      1 motorändplatta
      2 motorändplattan
      1 motorbanor
      1 motorbränsle
      1 motorbroms
      1 motorcortex
      1 motorcortexstimulering
      1 motorcykel
      1 motorcykelhjälm
      1 motorcykelsport
      6 motorer
      9 motorik
      2 motoriken
      1 motorikövningar
     20 motorisk
     38 motoriska
      4 motoriskt
      1 motorkomplex
      1 motorljudet
      2 motorn
      1 motornerver
      2 motorneuron
      1 motorneuronen
      2 motorneuronskada
      2 motorpackningar
      1 motorsignalering
      1 motorsvar
      1 motortrafikleder
      2 motorväg
      1 motorvagnståg
      2 motöverföring
      8 möts
      1 motsägande
      1 motsägelse
      2 motsägelsefull
      3 motsägelsefulla
      2 motsaten
     22 motsats
     29 motsatsen
      3 motsatser
     21 motsatt
     20 motsatta
      3 motsätter
      3 motsättning
      2 motsättningar
      1 motspelare
      5 motstå
     13 motstånd
      9 motståndare
      2 motståndaren
      1 motståndargrupperingarna
      1 motståndarna
      5 motståndet
      6 motståndskraft
      3 motståndskraften
      3 motståndskraftig
      4 motståndskraftiga
      1 motståndsresurser
      1 motsträviga
      5 motstridiga
      1 motstridigheter
      1 motströms
      3 motsvara
      3 motsvarade
     71 motsvarande
     43 motsvarar
      4 motsvaras
      1 motsvarat
      5 motsvarighet
      6 motsvarigheten
      2 motsvarigheter
      1 motsvarigheterna
      1 mött
      1 motta
      1 mottaga
      4 mottagande
      1 mottagarbakterien
      1 mottagarbakteriens
      3 mottagarcellen
      9 mottagare
      7 mottagaren
      6 mottagarens
      1 mottagarländer
      1 mottagarna
      1 mottagarorganismen
      1 mottagceller
      2 mottagit
      1 mottagits
      4 mottaglig
      9 mottagliga
      1 mottagligen
      5 mottaglighet
      3 mottagligheten
      1 mottagligt
      5 mottagning
      2 mottagningar
      1 mottagningarna
      1 mottagningen
      1 mottagrens
      5 mottar
      2 mötte
      4 möttes
      1 mottitaktiken
      1 motto
      1 mötts
      1 moturs
     37 motverka
      1 motverkan
     24 motverkar
      6 motverkas
      2 motvilja
      1 motvilligt
      1 motvisar
      1 mouches
      1 moulin
      2 mountain
      2 mounted
      1 mounting
      1 mouse
      1 move
      4 movement
      1 movementsömn
      1 mozart
      1 mozarteffekten
      1 mozarts
      1 mpa
      1 mpformat
      2 mpr
      6 mprvaccin
      1 mprvaccination
      5 mprvaccinet
      5 mpspelare
      8 mr
      1 mra
      1 mrbildtagning
      1 mrbildtagningstekniker
      1 mrbröst
      1 mrem
      2 mri
      1 mrimagnetic
      1 mristudier
     15 mrkh
      1 mrkhsyndromet
      4 mrna
      1 mrnatranskript
      1 mromänniskorätt
     16 mrsa
      1 mrsabakterier
      1 mrsabärare
      1 mrsainfektioner
      2 mrsastammar
      1 mrskanning
      7 mrt
      1 mrtsnittbild
     10 ms
      2 mscdsc
      1 mslt
      1 msm
      8 msv
      1 m�ta
      1 mtc
      1 mto
      1 mtuberculosis
      1 mtvgenerationen
      1 mtyp
      1 mucc
      1 mucin
      1 mucoangin
      1 mucosa
      1 [mucosa]
      2 mucosalagret
      1 muddring
      1 mukokutan
      3 mukösa
      1 muköst
      1 mul
      1 mula
      1 muladhara
      1 muldoon
      1 mulitelektroder
      1 mulkak
      1 mullard
      1 mullbärsväxter
      2 müller
      2 müllerian
      1 mülleriskt
      1 müllersk
      2 müllerska
      2 mülleruri
      1 mullrande
      1 mullvadssalamandrar
      1 multiaxial
      1 multiaxiala
      3 multibacillär
      1 multibegåvningen
      1 multicellulär
      1 multicenterstudie
      1 multiceps
      3 multidesign
      1 multidisciplinär
      1 multidisciplinära
      1 multielektrod
      1 multifaktorell
      1 multifaktorella
      2 multifaktoriell
      1 multifokal
      1 multiforme
      2 multilocularis
      1 multimedia
      2 multimeter
      2 multimetern
     11 multimetrar
      1 multimetrarna
      1 multimiljonmarknad
      1 multimodalt
      2 multinationella
      3 multinationellt
      1 multiorgandysfunktion
      2 multiorgansvikt
     11 multipel
      8 multipla
      1 multiplaflertal
      2 multiplanar
      1 multiplar
      1 multiple
      4 multiplicera
      1 multiplicerad
      1 multiplicerades
      1 multipliceras
      1 multiplicerat
      1 multiplied
      2 multipotenta
      1 multiproblemklienter
      1 multireceptiva
      6 multiresistent
      7 multiresistenta
      1 multiterapi
      1 multitrauma
      3 multivitamintabletter
      1 multocida
      1 mum
      1 mumie
      1 mumier
      1 mumiers
      1 mumifierade
      1 mumifieras
      1 mumla
      1 mumlande
     37 mun
      2 munarmar
      1 munbottnen
      1 muncancer
      1 munch
      1 münchen
      1 mundebo
      6 mundelar
      2 mundelarna
      1 mundiprincipen
      1 munduk
      1 mundusch
      1 munfull
     10 munhåla
     43 munhålan
      4 munhålans
      1 munhålecancer
      1 munhälsa
      1 munhälsan
      4 munhygien
      1 munhygienist
      2 munk
      7 munkar
      2 munkarna
      2 munken
      1 munkhatt
      1 munkmössa
      1 munmetoden
      1 munmotmunmetoden
      2 munnar
      1 munnäsa
     86 munnen
      6 munnens
      1 munnfull
      1 munöppning
      1 munöppningen
      1 munsår
      1 munsjukdomar
      1 munskador
      6 munskölj
      1 munsköljningar
      1 munskydd
      1 munslemhinnan
      2 munsönderfallande
      3 munspray
      1 munsprayer
      4 munstycke
      2 munstycket
      2 munsvalget
      2 muntligt
      8 muntorrhet
      1 munvård
      1 munvårdsprodukter
     14 munvatten
      1 munvattnet
      1 munverktygen
      3 mupirocin
      1 mur
      3 murad
      1 murar
      2 murarna
      1 murbinka
      3 murcs
      1 murcslikanande
      1 murcsliknande
      1 murder
      2 murphy
      1 murphys
      4 murray
      1 murrumbidgee
      1 murverk
      3 mus
      6 musarm
      1 musarmsbesvär
      1 musbett
      1 muscimol
      8 musculus
      1 muse
      1 musée
      2 museer
      1 museet
      1 musen
      8 museum
      1 mushrooms
     29 musik
      1 musikakupunktur
      1 musikalisk
      4 musikaliska
      1 musikaliskreligiösa
      1 musikaliskt
      6 musiken
      1 musikens
      4 musiker
      1 musikgrupper
      1 musikhögskolan
      4 musikinstrument
      1 musikkassett
      1 musiks
      3 musikstycke
      1 musikstycken
      1 musikterapeut
      2 musikterapeuter
      1 musikterapeutiska
      6 musikterapi
      1 musikterapier
      1 musiktraditionen
      1 musikupplevelse
      1 musikverk
      1 muskarin
      2 muskarinerga
      2 muskarinreceptorer
      3 muskarinreceptorerna
     27 muskel
      2 muskelaktivitet
      1 muskelanspänning
      2 muskelarbete
      3 muskelatrofi
      1 muskelavslappande
      2 muskelavslappnande
      1 muskelavslappning
      1 muskelbädd
      1 muskelband
      3 muskelbiopsi
      8 muskelbristning
      1 muskelbristningar
      2 muskelbyggare
      4 muskelcell
      1 muskelcellen
      3 muskelceller
      8 muskelcellerna
      1 muskeldomningar
      2 muskeldystrofi
      1 muskeldystrofier
      1 muskelfack
      1 muskelfackens
      1 muskelfascikel
      5 muskelfästen
      4 muskelfiber
      2 muskelfibrer
      1 muskelförändringar
      1 muskelförlamning
      2 muskelförtvining
      1 muskelfunktion
      1 muskelgenererad
      1 muskelgrupp
      2 muskelgrupper
      1 muskelinflammation
      2 muskelknutar
      4 muskelknutor
      2 muskelkontraktion
      1 muskelkontrollen
      1 muskelkoordination
      2 muskelkraft
      1 muskelkraften
      2 muskelkramper
      1 muskellager
     12 muskelmassa
      1 muskelmassan
     38 muskeln
      3 muskelns
      1 muskelorgan
      1 muskelprestation
      1 muskelproteiner
      1 muskelprov
      1 muskelretning
      1 muskelreumatism
      5 muskelrörelser
      1 muskelryckningar
      1 muskelsammandragning
      4 muskelsammandragningar
      1 muskelsinne
      1 muskelsinnet
      3 muskelsjukdom
      1 muskelsjukdomar
      2 muskelskada
      1 muskelskador
      1 muskelskeletala
      2 muskel�skelettskador
      1 muskelskida
      1 muskelskikt
      3 muskelsmärta
      5 muskelsmärtor
      1 muskelsmärtorna
      1 muskelsönderfall
      3 muskelspänning
      3 muskelspänningar
      1 muskelspasm
      1 muskelspasmer
      1 muskelspolarna
      2 muskelstelhet
      1 muskelstorleken
      1 muskelsträckning
      4 muskelstyrka
      2 muskelstyrkan
     12 muskelsvaghet
      1 muskelsymtom
      1 muskeltillväxt
      8 muskeltonus
      1 muskeltonusen
      1 muskeltonusförlust
      2 muskelträning
      1 muskeltrauman
      2 muskeltrötthet
      1 muskeluppbyggnaden
      1 muskelvägg
      1 muskelväggar
     19 muskelvärk
      7 muskelvävnad
      2 muskelvävnaden
      1 muskelvolymökning
     81 muskler
     70 musklerna
      2 musklernas
      1 muskotnötter
      3 muskulär
      5 muskulära
      2 muskulärt
     24 muskulatur
     15 muskulaturen
      1 muskulaturens
      3 muskuloskeletala
      4 muslimer
      1 muslimsk
      9 muslimska
      2 musselsäsongen
      1 musseroner
      1 musseronerna
      1 musslor
      1 musstam
      1 mutans
      1 mutanter
     39 mutation
     12 mutationen
     29 mutationer
      2 mutationerna
      1 mutationsom
      1 mutationsrisk
      3 mutera
      2 muterad
      2 muterade
      1 muteras
      1 muterat
     17 mutism
      1 mutismen
      1 mutistisk
      1 mutsuru
      1 mutter
      1 mutterkreuz
      1 mutualism
      1 mutus
      9 mv
      1 �mv
      1 mva
      2 mvaa
      1 mvab
      1 mwl
      1 mwt
      3 myalgi
      1 myastena
      1 myasthenia
      5 mycel
      1 mycelet
      1 mycelieliknande
      1 myceliemassa
      1 myceliemassans
      1 mycelievävnad
      1 mycelsträngar
      2 mycin
      1 mycken
   1123 mycket
      1 mycobacteriaceae
     14 mycobacterium
      1 mycoidesorganism
      3 mycoplasma
      2 mydriasis
      1 mydriatriska
      1 mydrostatikum
      3 myelin
      3 myelinet
      1 myeliniserat
      2 myelinolys
      1 myelinprojektet
      2 myelit
      1 myeloblast
      1 myelocyt
      1 myelogent
      2 myeloid
      3 myeloisk
     14 myelom
      1 myelomcell
      1 myelomcellen
      3 myelomeningocele
      1 myelomet
      1 myelomskelett
      1 myelopati
      5 mygg
      2 mygga
     11 myggan
      1 myggangrepp
      4 myggans
      2 myggart
      1 myggarter
      1 myggbeståndet
      8 myggbett
      5 mygglarver
      5 myggmedel
      3 myggnät
     13 myggor
      3 myggorna
      1 myggornas
      1 myggplåga
      1 myggpopulationerna
      1 myggstammarna
      3 myggstick
      1 myhos
      1 myhrman
      1 mykobacterium
      1 mykobakteriell
      1 mykobakterieproteiner
      6 mykobakterier
      2 mykobakterierna
      1 mykocerosinsyror
      2 mykolsyra
      1 mykoöstrogener
      2 mykoplasma
      1 mykoplasmainfektion
      1 mykoplasmainfektioner
      2 mykorrhiza
      1 mylan
      1 mylla
      9 myndig
      9 myndiga
     18 myndighet
     14 myndigheten
      2 myndighetens
     24 myndigheter
     11 myndigheterna
      1 myndigheternas
      2 myndigheters
      5 myndighetsålder
      2 myndighetsåldern
      1 myndighetskontroll
      1 myndighetsuppgifter
      1 mynna
     18 mynnar
      5 mynning
      1 mynningen
      5 mynt
      1 mynta
      7 myntade
     24 myntades
      3 myntat
      1 myntats
      1 myntrullebildning
      1 myntrullebildningen
      1 myo
      1 myocardium
      1 myocardskintigrafi
      1 myodes
      1 myoelasticitet
      1 myoepitelceller
      1 myoepitelcellerna
      3 myoglobin
      5 myokardiet
      5 myokardit
      3 myokardium
      1 myokloni
     34 myom
      1 myomen
      1 myomens
      8 myomet
      1 myometriet
      1 myometrisk
      1 myometrium
      1 myomets
      1 myomtumörer
      1 myonycteris
      3 myopati
      1 myopatisk
      1 myos
      3 myosit
      4 myostatin
      1 myostatinhämmare
      1 myoview
      1 myr
      1 myra
      1 myrar
      2 myrberg
      1 myrdaling
      2 myrkrypningar
      4 myror
      1 myrpiggsvin
      1 myrra
      1 myrraolja
      1 myrstackar
      4 myrsyra
      1 myrsyrans
      1 mysterier
      1 mysteriska
      2 mysterium
      1 mysticism
      3 mystik
      1 mystiken
      3 mystiker
      1 mystiska
      4 myt
      1 mytbildningen
      9 myten
      4 myter
      1 myterna
      3 myth
      1 mytisk
      1 mytiska
      6 mytologi
      1 mytologier
      7 mytologin
      1 mytologiserad
      1 mytologiska
      1 mytoman
      2 mytomanen
      2 mytomaner
      3 mytomani
      1 mytomanin
      1 mytomans
      4 myxödem
      4 myxom
      2 myxomet
     26 n
      4 na
     59 nå
      1 naafa
      1 naaq
      4 näbb
      1 �näbb
      1 näbbdjur
      4 näbben
      1 näbbens
      2 näbbliknande
      1 näbbmöss
      1 nacclhco
      1 nacetylmetoxitryptamin
      1 nacfhco
      1 nachtmahr
      1 nachtmerrie
      2 nack
      1 nackbehandlingar
      1 nackbenets
      3 nackbesvär
      6 nackdel
     13 nackdelar
      4 nackdelarna
      8 nackdelen
     13 nacke
     21 nacken
      1 nackens
      1 nackkrage
      1 nackmanipulation
      1 nackområdet
      1 nackrelaterad
      1 nackskada
      1 nackskuldersmärta
      2 nacksmärta
      1 nacksmärtor
      3 nackspärr
      1 nackstelhet
      1 nackstöd
      3 nackstyvhet
      1 nackvävnad
      3 nacl
      1 nacllösning
      3 naclo
      1 nacls
      1 nacn
      1 nad
     19 nådde
      1 nåddes
      1 nadh
      1 nadhberoende
      3 nadi
      1 nadier
      1 naevi
      1 naevocellulära
      1 naevus
      2 naf
      5 naftalen
      1 naftol
      1 nagana
      1 någe
      3 nagel
      1 nagelangrepp
      1 nagelbädden
      2 nagelbitning
      1 nagelemalj
      1 nagelemaljen
      2 nagelfil
      3 nagelfilar
      1 nagelfilning
      1 nagelkanten
      5 nagelklippare
     10 nagellack
      2 nagellacket
      1 nagellacksborttagare
      2 nageln
      1 nagelns
      1 nagelpetare
      1 nagelproblem
      1 nagelsjukdomar
      1 nagelsvamp
      1 nageltång
      2 nageltrång
     11 naglar
      8 naglarna
      1 nagna
    593 någon
      1 någondera
      1 någonnågra
      1 någons
      6 någonsin
      7 någonstans
     16 någonting
      9 någorlunda
    521 något
      2 någotsånär
    478 några
      1 nahco
      2 nahuatl
      2 nai
      1 naivitet
      1 nåjd
      2 nåjden
      1 najonerna
      1 najonkanaler
      1 nakanaler
      1 nakazono
      2 naken
      2 nakenbad
      3 nakenhet
      1 nakenyoga
      5 nakna
      1 nakpumpen
     21 nål
     13 nålar
      2 nålarna
      1 nålbiopsi
      1 nåldelning
      1 nålelektrod
      1 nålelektroder
      2 nålelektromyografi
      3 nålen
      1 nålens
      1 nålformiga
      2 nålfri
      1 nålinstrument
      1 naloxon
      2 nålstick
      3 nålsticken
      1 nålstickens
      1 nålsticket
      1 nålsticksretningen
      1 namedevelop
      1 namelobotomidanmark]
      1 nament
      1 namewwwcdcgovparasitestrichinellosis
      1 namewwwsmittskyddsinstitutetsesjukdomartrikinos
      1 namewwwsvasesvdjurhalsazoonosertrikinossomzoonos
      1 namikoshi
     42 nämligen
    145 namn
      3 nämna
      1 nämnande
      1 nämnare
      3 nämnaren
     27 nämnas
      1 namnbytet
      1 namnceremonier
      3 nämnd
     21 nämnda
      1 nämnde
      2 nämnden
      3 nämnder
      1 nämnderna
      1 nämnders
      4 nämndes
     11 namnen
      6 nämner
    219 namnet
      2 namnets
      4 namnformer
      1 namnformerna
      1 namnförslag
      3 namngav
      2 namngavs
      3 namnge
      1 namnger
      4 namnges
      1 namngett
      1 namngiven
      2 namngivet
      2 namngivna
      2 namngivning
      1 namngivningen
      1 namnkunnigaste
      1 namnlika
      1 namno
     11 nämns
      1 namnsorter
      4 nämnt
      2 nämnts
      3 nämnvärd
      1 namnvarianter
      5 nämnvärt
      1 nampulaprovinsen
      1 nana
      2 nancy
      1 nano
      1 nanogram
      2 nanomaterial
      4 nanometer
      1 nanopartiklar
      1 nanopartiklarna
      1 nanosekund
      1 nanosekunder
      1 nanoteknologi
      3 naoh
      1 napi
      4 napoleon
      3 napoleonkrigen
      1 napoleons
      1 napoleonsk
      2 nappflaskor
      2 naprapat
      1 naprapaten
      7 naprapater
      1 naprapaterna
      1 naprapatförbundet
      1 naprapathic
      1 naprapathögskolan
      1 naprapathögskolanär
      5 naprapati
      1 naprapatin
      1 naprapatins
      1 naprapatutbildning
      1 naprapatutbildningarna
      1 naprapatutbildningen
      1 napravit
      2 naproxen
     67 når
   1330 när
    144 nära
      1 näradöden
      2 näradödenupplevelse
      3 näradödenupplevelser
      4 näraliggande
      1 närapå
      1 närbeläget
      1 närbesläktad
      8 närbesläktade
      4 närbesläktat
      1 närbutik
      1 narciss
      2 narcisser
      1 narcisserna
     10 narcissism
      2 narcissisten
      5 narcissistisk
      1 narcissläktet
      1 narcissläktets
      3 narcissus
      1 narcotic
      1 narcotics
      1 närde
      1 närhelst
      9 närhet
     36 närheten
      1 närhets
      1 närhetssökande
     26 näring
      4 näringen
      1 närings
      5 näringsämne
     31 näringsämnen
      3 näringsämnena
      1 näringsbalansen
      4 näringsbehov
      1 näringsberäkning
      1 näringsberäkningar
     13 näringsbrist
      1 näringsceller
      1 näringsfaktorer
      1 näringsförlust
      1 näringsförlusten
      2 näringsförluster
      1 näringsfysiologi
      1 näringsgrenar
      1 näringsidkare
      2 näringsinnehåll
      1 näringsintag
      3 näringsintaget
      1 näringskällan
      4 näringskedjan
      9 näringslära
      3 näringsliv
      1 näringslivet
      4 näringslösningar
      1 näringsmässig
      1 näringsmässigt
      1 näringsmineraler
      4 näringsrik
      2 näringsrika
      3 näringsriktig
      2 näringsrubbning
      5 näringsrubbningar
      1 näringsstatus
      6 näringstillförsel
      2 näringstillgång
      1 näringstillskott
      1 näringstillståndet
      5 näringsupptag
      1 näringsupptagandet
      2 näringsupptaget
      1 näringsvärde
      1 näringsvärdet
      1 närinställning
      2 narke
      1 närke
      1 narkissos
     33 narkolepsi
      1 narkolepsifall
      1 narkolepsifallen
      1 narkolepsiforskning
      3 narkoleptiker
      1 narkoman
      1 narkomanen
      9 narkomaner
      1 narkomanerna
     11 narkomani
      1 narkomaniepidemi
      1 narkomanvård
      4 närkontakt
     40 narkos
      1 narkosdjup
      1 narkosdjupet
      2 narkosläkare
      1 narkosläkaren
      5 narkosmedel
      1 narkosmedlen
      1 narkosmedlet
      1 narkosmetoden
      2 narkospersonalen
      1 narkosrelaterade
      1 narkotik
     39 narkotika
      1 narkotikaanvändning
      1 narkotikaavvänjning
      1 narkotikaberoende
      2 narkotikabrott
      1 narkotikabrottskonvention
      1 narkotikabrottskonventionen
      1 narkotikabrottslighet
      1 narkotikabrottsling
      1 narkotikadebatten
      1 narkotikaförgiftning
      2 narkotikafria
      2 narkotikafritt
      1 narkotikahanteringen
      9 narkotikaklassad
      5 narkotikaklassade
      3 narkotikaklassat
      1 narkotikaklassats
      2 narkotikakonsumtion
      2 narkotikakonvention
      3 narkotikakonventioner
      1 narkotikalagstiftningen
      1 narkotikamarknaden
      2 narkotikamissbruk
      2 narkotikamissbrukare
      1 narkotikan
      1 narkotikans
      1 narkotikaområdet
      6 narkotikapolitik
      2 narkotikapolitiken
      1 narkotikapolitisk
      1 narkotikarelaterade
      1 narkotikaupplysning
      4 narkotisk
      4 narkotiska
     12 närliggande
      6 närma
      1 närmade
      7 närmar
     40 närmare
     25 närmast
     25 närmaste
      1 närmat
      2 närmiljö
      1 närmiljön
      2 närminnet
      3 närmre
      1 närpolisen
      1 närproducerat
      2 närpunkten
      1 närsalter
      1 närsalterna
      1 närseendets
      1 närsläktade
     15 närstående
      1 närståendei
      1 närståendes
      1 närstridsvapen
      1 närsynt
      1 närsynta
      5 närsynthet
      1 närsynthetsutvecklingen
      1 narus
      3 närvara
     49 närvarande
     24 närvaro
      8 närvaron
      1 �närvaron
      1 närvaroövningar
      3 nås
      2 näs
     48 näsa
      1 nasal
      1 nasala
      1 nasalt
     65 näsan
      1 näsanär
      9 näsans
      1 näsaöronpassagen
      2 näsbenet
      6 näsblod
      3 näsblödning
      4 näsblödningar
      1 näsblödningen
      4 näsborrar
      6 näsborrarna
      1 näsborrarnas
      2 näsborre
      4 näsborren
      1 näsbryggan
      1 näsbryggor
      3 näsdroppar
      4 näsduk
      5 näsdukar
      8 näsduken
      1 näsduksväska
      1 näsepitlet
      1 näsgången
      1 näsgrimma
      2 näshåla
     12 näshålan
      1 nasitergium
      1 näsläppveck
      2 näslund
      1 näsmask
      1 naso
      1 nasofaryngit
      2 nasofarynx
      3 nasogastrisk
      1 nasonex
      2 näsöppningarna
      2 näsor
      4 näspetande
      2 näspetning
      2 näspiercing
      4 näspiercingar
      1 näspiercingarna
      2 näspiercingen
      4 näsplastik
      1 näsprov
      1 näsring
      1 näsroten
      2 näsryggen
      1 nässelcell
      6 nässelceller
      5 nässelcellerna
     12 nässeldjur
      4 nässeldjuren
      2 nässeldjurens
      1 nässeldjurskolonier
      1 nässelduk
      2 nässelfeber
      1 nässelfibrerna
      1 nässelfjäril
      1 nässelkål
      1 nässelkapslar
      2 nässelsläktet
      1 nässelsnärja
      1 nässelsoppa
      1 nässelstånd
      3 nässelutslag
      1 nässelvatten
      1 nässelväxter
      2 nässköljning
      1 nässköljningkanna
      1 nässköljningskannan
      1 nässla
      2 nässlem
      3 nässlemhinnan
      1 nässlor
      1 nässlorna
      1 nässmycket
      1 nässpolning
      3 nässpray
      1 nässprayer
      3 nässprej
      1 nässprejer
      1 nässtyng
      1 nässtyngfluga
      3 nässvalget
     26 näst
     45 nästa
    180 nästan
     10 nästäppa
      2 nästintill
      1 nästippar
      2 nästkommande
      1 nästlar
      1 nästorkare
      1 näsvidgare
      2 näsvinge
      1 näsvingevidgare
      1 nat
      5 nät
      3 natalensis
      1 nätbur
      1 nätbutik
      1 nätbutikerna
      2 nätet
      1 nätfrånkopplare
      1 nathan
      3 näthandeln
      1 näthandlare
      1 näthandlarna
      4 näthinna
     13 näthinnan
      6 näthinneavlossning
     26 national
      1 nationalblomma
      3 nationale
      1 nationalekonomin
      2 nationalencyklopedin
      1 nationalitetsmärke
      1 nationalkaraktären
      4 nationalpark
      1 nationalreligion
      9 nationell
     29 nationella
      3 nationellt
      2 nationen
      1 nationer
      5 nationerna
      2 nationernas
      2 nations
      3 nativa
      2 nativitet
      1 nätmagen
     16 natrium
      1 natriumacetoacetat
      1 natriumalginat
      1 natriumatomer
      1 natriumbalans
      5 natriumbensoat
      2 natriumbikarbonat
      1 natriumcyanid
      1 natriumdodecylsulfat
      1 natriumfenolat
      6 natriumfluoracetat
      2 natriumfluorid
      2 natriumföreningen
      1 natriumhalterna
     12 natriumhydroxid
      1 natriumhydroxidlösning
     10 natriumhypoklorit
      8 natriumjoner
      1 natriumjonerna
      1 natriumkanalblockering
      1 natriumkarbonat
      1 natriumkloracetat
      1 natriumklorat
     15 natriumklorid
      1 natriumkloridlösning
      1 natriumklorit
      2 natriumkromoglikat
      1 natriumlauryletersulfat
      2 natriumlaurylsulfat
      1 natriumnitrat
      2 natriumnitrit
      1 natriumpermanganat
      1 natriumpumpar
      4 natriumsalt
      2 natriumsalter
      3 natriumsulfat
      1 natriumtvål
      1 natriumtvålar
      1 natriumvalproat
      1 natriuretisk
      2 natriuretiska
      3 natronlut
      1 nätspänning
     13 natt
     25 nått
      3 nattaktiv
      1 nattbindor
      4 nattblindhet
      2 nattblöja
      1 nattblöjor
      1 nättelduk
     42 natten
      2 nattens
      7 nätterna
     14 nattetid
      1 nattfjärilen
      1 nattflygningar
      1 natthosta
      1 nättidning
      4 nattklubbar
      2 nattkorsetter
      1 nattkylan
      1 nattläger
      4 nattlig
      9 nattliga
      1 nattligt
      1 nattmänniska
      1 nattöppna
      3 natts
      1 nattskategräs
      4 nattskatta
      2 nattskattan
      6 nattskräck
      5 nattsömn
      1 nattsömnen
      1 nattvardsgåvorna
     25 natur
      1 naturae
      1 natural
      3 naturalförlopp
      4 naturalförloppet
      3 naturaliserad
      1 naturaliserade
      1 naturaliserats
      1 naturalistisk
      1 naturande
      2 naturbehov
      1 naturbetesmark
      1 naturborstar
      4 nature
     41 naturen
      1 naturenbakom
      5 naturens
      1 naturfiber
      1 naturfibrer
      1 naturfibrerna
      1 naturfilosof
      1 naturfilosofi
      1 naturfilosofin
      1 naturfilosofiska
      4 naturfolk
      1 naturfolks
      2 naturgas
      1 naturgummi
      1 naturhår
      1 naturhistoria
      1 naturistkretsar
      1 naturkatastrof
      6 naturkatastrofer
      2 naturläkemedel
     27 naturlig
     65 naturliga
      2 naturligaste
      1 naturligen
     85 naturligt
      7 naturligtvis
      2 naturmaterial
      1 naturmedel
      1 naturmediciner
      1 naturopaten
      1 naturrätten
      2 naturreservat
      1 naturskyddsföreningen
      1 natursten
      1 natursvamp
      1 naturtampong
      1 naturtrogna
      2 naturvårdsunionen
      1 naturvårdsunionens
      1 naturvårdsverket
      1 naturvetarna
      4 naturvetenskap
      1 naturvetenskapens
      2 naturvetenskapliga
      1 naturvetenskapligt
     25 nätverk
      9 nätverket
      2 nätverkets
      1 nätverksanalysator
      2 nätverksanalysatorer
      2 nätverksparametrar
      1 nauru
      1 nav
      1 navel
      1 navelartärvenkateter
      2 navelbråck
      2 navelhöjd
     13 naveln
      1 navelpiercingar
      4 navelsträngen
      1 näver
      2 navigering
      1 navlad
      1 navlar
      1 nazaret
      3 nazareto
      1 nazismens
      1 nazist
      1 nazisten
      1 nazister
      3 nazisternas
      1 nazistisk
      3 nazistiska
      8 nazityskland
      1 nazitysklands
      1 nbc
      1 nbedelefolkets
      1 nbn
      1 nca
      2 ndd
      1 ndealkylation
      1 ndes
      1 ndm
      2 ne
      2 neapel
      1 neapolitanska
      1 neardeath
      1 neardeathexperiences
      1 neas
      2 nebulisator
      1 nécessaire
      1 necessär
      1 necessären
    105 ned
     52 nedan
     16 nedanför
      9 nedanstående
      1 nedärvas
      1 nedärvd
      3 nedärvda
      1 nedärvs
      1 nedärvt
     14 nedåt
      1 nedåtflytande
      1 nedåtgående
      2 nedåtriktad
      1 nedåtriktade
      1 nedåtrullade
      1 nedbringade
      1 nedbruten
      1 nedbrutet
      1 nedbrutna
      6 nedbrytande
      1 nedbrytbara
      1 nedbrytbart
      1 nedbryter
     36 nedbrytning
     10 nedbrytningen
      1 nedbrytningsämnen
      1 nedbrytningsprocess
      2 nedbrytningsprocesser
      4 nedbrytningsprodukt
      5 nedbrytningsprodukter
      1 nedbrytningsreaktioner
      2 nederbörd
      1 nederdel
      1 nederkanten
      1 nederlaget
      1 nederländaren
      1 nederländarna
     26 nederländerna
      1 nederländernas
      2 nederländsk
      3 nederländska
      6 nedersta
      2 nedför
      2 nedförsbacke
      1 nedförslut
      5 nedfrysning
      1 nedfrysnings
      3 nedgång
      1 nedkyld
      9 nedkylning
      1 nedkylningen
      1 nedladdning
      1 nedlagda
      1 nedläggas
      1 nedlägges
      1 nedläggning
      1 nedlåtande
      1 nedliggande
      2 nedlöpande
      1 nedmontering
      1 nedokromil
      1 nedom
      1 nedprioriteras
     84 nedre
      1 nedreglerar
      2 nedsänkt
    121 nedsatt
      5 nedsatta
      5 nedsättande
      3 nedsätter
     17 nedsättning
      7 nedsättningar
      1 nedsättningarna
      2 nedsätts
      1 nedskrivet
      1 nedskrivna
      1 nedsläckt
      1 nedslående
      1 nedslag
      1 nedsliten
      1 nedslitet
      1 nedslitna
      1 nedslitningsprocessen
      1 nedsmittade
      1 nedsmutsad
      2 nedsövd
      1 nedsövning
      2 nedstämd
      1 nedstämda
      7 nedstämdhet
      2 nedstämdheten
      1 nedstämt
      2 nedstigning
      2 nedströms
      1 nedsvalda
      1 nedsväljning
      1 nedtecknad
      1 nedtecknade
      1 nedtecknades
      1 nedtecknande
      1 nedtill
      1 nedtittande
      1 nedträngda
      1 nedtryckt
      1 nedtryckthet
      1 nedvandring
      1 nedvärdera
      1 nedvärderande
      1 needs
      1 neelix
      1 neet
      1 nefadar
      6 nefazodon
      2 nefrektomi
      1 nefridier
      2 nefrit
      1 nefrologi
      3 nefropati
      2 nefrotiskt
      1 negation
     32 negativ
    105 negativa
      2 negative
      1 negativism
      2 negativistiskt
     48 negativt
      1 negev
     16 neglect
      1 neglected
      1 neglekt
      1 neglektalexi
      1 nei
      1 neil
      1 neinstein
     12 neisseria
      4 nej
      1 nejfråga
      1 nejlikeolja
      2 nejlikväxter
      4 neka
      2 nekades
      3 nekande
      1 nekas
      1 nekat
      1 nekats
     14 nekros
      1 nekrotiserad
      2 nekrotiserande
      2 nekrotiska
      4 nektar
      1 nektarier
      1 nélaton
      1 nematocera
      1 nematocyster
      1 nematocyter
      1 nematocyterna
      2 nematoda
      1 nematoder
      1 nematoderna
      7 nemg
      1 nemgundersökningen
      2 nemorosa
      1 neocortex
      2 neoformans
      3 neokortikala
      3 neolitikum
      1 neolitisk
      1 neologism
      2 neologismer
      1 neonatal
      1 neonatalavdelning
      1 neonatalavdelningen
      1 neonatalvård
      1 neonatalvården
      1 neonatologer
      1 neonatorum
      1 neonatus
      9 neoplasi
      1 neoplasier
      3 neoplastisk
      1 neorganics
      1 neosalvarsan
      1 neosalvarsanet
      1 neoten
      1 neovitalism
      1 nepal
      2 nephropathia
      1 neptunigördel
    257 ner
      6 neråt
      7 nere
      1 nerfläckning
      4 nerium
      1 nerkonverteras
      1 nerkylning
      1 nermalda
      3 nerman
      1 nermans
      1 nero
      1 nersmältning
      3 nertill
      5 nerv
      1 nervaktionspotentialerna
      1 nervaktivitet
      2 nervändar
      1 nervände
      1 nervänden
      1 nervändplattans
      2 nervändsluten
      1 nervändslutet
      4 nervbanor
      3 nervbanorna
      1 nervblockad
     13 nervcell
     10 nervcellen
      5 nervcellens
     47 nervceller
      8 nervcellerna
      2 nervcellers
      1 nervcells
      1 nervcellsdöd
      1 nervcellsnybildningen
      1 nervcellstillväxt
      1 nervcellsutskott
      1 nervcentra
      1 nervdiket
      1 nerve
      1 nerveller
      6 nerven
     42 nerver
     10 nerverna
      5 nervernas
      1 nervfeber
      1 nervfiber
      1 nervfibererna
      1 nervfiberlager
      3 nervfibrer
      1 nervgas
      1 nervgaser
      1 nervgaserna
      3 nervgift
      1 nervig
      2 nervimpuls
      1 nervimpulsen
      1 nervimpulsens
     14 nervimpulser
      1 nervinflammationer
      2 nervinklämning
      2 nervkanalen
      1 nervknippen
      1 nervknutor
      1 nervledningshastigheten
      1 nervledningsundersökningar
      2 nervmuskelsjukdomar
      1 nervnäringsmedlet
      1 nervnät
      3 nervös
     22 nervosa
      2 nervösa
      7 nervositet
      2 nervpåverkan
      1 nervprojektioner
      1 nervprojektionerna
      2 nervrötter
      1 nervryckningar
      1 nervs
      2 nervsignaler
      1 nervsignalerna
      2 nervsjukdomar
      4 nervskada
      6 nervskador
      7 nervsmärta
      1 nervsmärtor
      2 nervssystemet
      3 nervstimulering
      1 nervstimulus
      1 nervsvaghet
      7 nervsystem
    175 nervsystemet
      8 nervsystemets
      1 nervsystems
      1 nervsytemet
      1 nervterminaler
      3 nervtillväxtfaktor
      1 nervtråd
      1 nervtrådar
      1 nervtråden
      1 nervtrådskapseln
      9 nervus
      4 nervvävnad
      1 nes
      1 nested
      1 nestlé
      2 netherlands
      1 nettoflöde
      2 nettokolhydrater
      1 nettoladdningen
      1 nettotillskott
      2 netzel
      1 neuhauser
      1 neumann
     12 neurala
      1 neuralfåran
      4 neuralgi
      2 neuralrör
      2 neuralröret
      2 neuraminidas
      1 neuraminidashämmare
      8 neurasteni
      1 neurit
      1 neuroanatomer
      2 neurobiologi
      1 neurobiologins
      1 neurobiologisk
      2 neurobiologiska
      3 neuroblastom
      1 neurobloc
      2 neuroborrelios
      1 neurochir
      4 neurodegeneration
      1 neurodegenerativ
      3 neurodegenerativa
      1 neurodegenerativt
      1 neurodiagnostisk
      1 neurodyni
     12 neuroendokrina
      4 neuroendokrinologi
      2 neuroendokrinologin
      1 neuroendokrinologiska
      1 neuroendokrinologiskt
      1 neuroetologi
      1 neurofibrom
      6 neurofibromatos
      1 neurofibromen
      1 neuroforskare
      1 neurofysiologen
      6 neurofysiologi
      2 neurofysiologisk
      2 neurofysiologiska
      1 neurogen
      2 neurogena
     32 neurogenes
      1 neurogenesberoende
      1 neurogenesen
      1 neurogeneshämmare
      1 neurogenområdena
      1 neuroglycopent
      2 neurografi
      3 neurohormoner
      9 neurohypofysen
      1 neuroimaging
      1 neuroimmunologiska
      2 neurointensivvård
      1 neurointensivvårdavdelning
      1 neurointensivvården
      1 neurokirugi
      2 neurokirurg
      2 neurokirurger
      1 neurokirurgerna
     12 neurokirurgi
     15 neurokirurgin
      2 neurokirurgins
      4 neurokirurgisk
     13 neurokirurgiska
      1 neurokirurgiskt
      1 neurokirurigiska
      1 neurokognitiv
      3 neurokognitiva
      1 neuroleptica
     16 neuroleptika
      1 neuroleptikabehandling
      1 neuroleptikabesläktade
      1 neuroleptikapreparat
      1 neuroleptikas
      3 neuroleptikasyndrom
      1 neuroleptikat
      6 neuroleptikum
      1 neuroleptikumläkemedel
      1 neuroleptiska
      1 neurolobus
      4 neurolog
      4 neurologen
      5 neurologer
      1 neurologerna
      3 neurologi
      3 neurologin
     31 neurologisk
     61 neurologiska
      7 neurologiskt
      1 neurology
      1 neuromodulator
      2 neuromuskulär
      4 neuromuskulära
      1 neuromuskulärt
     11 neuron
      3 neuronal
      5 neuronala
      2 neuronen
     11 neuroner
      6 neuronerna
      1 neuronernas
      1 neuroners
      4 neuronet
      1 neuronförlust
      1 neuronmigrationens
      1 neuronöverlevnad
      1 neuropati
      1 neuropatier
      3 neuropatisk
      1 neuropatologiska
      3 neuropeptid
      2 neuropeptider
      1 neuropeptiderna
      8 neuroplasticitet
      1 neuroplasticiteten
      1 neuroplasticitetens
      2 neuropsychiatric
      2 neuropsykiatri
      3 neuropsykiatrin
      7 neuropsykiatrisk
     12 neuropsykiatriska
      1 neuropsykiatriskt
      2 neuropsykologisk
      3 neuropsykologiska
      4 neuroradiologi
      1 neuroradiologin
     16 neuros
      1 neurosarkoidos
      2 neurosedyn
      1 neurosedynskadorna
      2 neurosedynskandalen
      1 neurosekretoriska
     25 neuroser
      3 neuroserna
      1 neurosfära
      1 neurosfärt
      1 neurosomatisk
      1 neurospecialiteter
      2 neurosphere
      1 neurosterapi
      7 neurosyfilis
      2 neuroticism
      5 neurotisk
      6 neurotiska
      3 neurotiskt
      2 neurotoxin
      1 neurotoxiskt
      5 neurotransmittor
      4 neurotransmittorer
      1 neurotransmittorerna
      3 neurotransmittorn
      1 neurotrofisk
      1 neurotropa
      1 neurotropiskt
      3 neurotyp
      1 neurotypa
      3 neurotypisk
      1 neurotypiska
      1 neurovaskulära
      2 neurovetenskap
      2 neurovetenskapen
      1 neurovetenskapliga
      3 neutral
      4 neutrala
      1 neutralisationstest
      4 neutralisera
      4 neutraliserar
      1 neutraliseras
      1 neutraliserat
      1 neutralisering
     10 neutralt
      3 neutrofila
      3 neutrofiler
      2 neutrofilerna
      7 neutroner
      1 neutronstrålning
      1 neutropeni
      1 nevada
      1 nevadensis
      1 never
      1 nevus
     35 new
      1 newage
      1 newcastle
      2 newcastlesjuka
      1 newdelhi
      1 newdelhimetallobetalaktamas
      1 newdelhimetallolaktamas
      1 news
      1 newtons
      1 nexus
      2 nez
     12 nf
      2 ngf
      2 ngkg
      1 ngl
      2 ngml
      1 ngn
      6 ngonorrhoeae
      2 ngonorrhoeaes
      4 nh
      1 nhk
      1 nhmrc
      1 nhs
      6 ni
      2 niacin
      1 niacinsyntesen
      1 niåver
      1 nice
      2 nicholson
      1 nicka
     16 nickel
      3 nickelallergi
      2 nickelallergiker
      1 nickeleksem
      1 nickelkadmiumackumulatorer
      1 nickelsilver
      1 nickeltitan
      1 nickeltitanlegering
      1 nicklet
      1 nicolae
      1 nicolas
      1 nicole
      1 nicolet
      1 nicot
      1 nicotiana
      1 nidana
      1 nidra
      1 niederschlesien
      1 niels
      1 nielsen
      2 nietzsche
      1 nifedipin
      1 nigella
      4 niger
      6 nigeria
      1 nightmare
      3 nigra
      2 nigricans
      1 nigrivalvis
      1 nigriventer
      1 nigrum
      2 nih
      1 nihilism
      1 nihilister
      1 nihl
      1 nihtredarna
      1 nikandros
      3 nikolaj
      1 nikon
      8 nikotin
      1 nikotinerg
      1 �nikotinerga
      1 nikotinersättning
      1 nikotinet
      1 nikotinkicken
      2 nikotinplåster
      1 nikotinreceptorer
      1 nikotintuggummi
      1 niktotinreceptorerna
      1 nile
      1 nileviruset
      4 nils
      5 nilsson
      1 nimh
      1 nina
      1 ninon
      1 nintendotumme
     30 nio
      1 niohundra
      1 nionde
      1 nioprocentregeln
      1 nipacide
      2 nipplegate
      1 nipponium
      2 nirvana
      1 nirvanasångaren
      1 nisal
      3 nisch
      2 nit
      1 nitbrillor
      1 nitbrillorna
      1 nitinol
      1 nitrat
      1 nitrater
      1 nitratet
      1 nitreras
      1 nitricum
      2 nitrobensen
      1 nitrobenzol
      3 nitrocellulosa
      4 nitrofurantoin
      2 nitroglycerin
      1 nitrohydroxifenylarsonsyra
      1 nitrosaminer
      1 nitrox
      1 nittio
      1 nittiotalet
      1 nittiotalismen
      2 nittonhundratalet
      1 niue
      1 niva
     82 nivå
      1 nivådiagnostik
     97 nivåer
     35 nivåerna
      1 nivåförändringarna
      1 nivalis
     18 nivån
      1 nivåpatogen
      1 nivåskillnader
      1 nivea
      1 nivens
      4 njur
     14 njurar
     53 njurarna
      4 njurarnas
      1 njurartärernas
      2 njurbäckenet
      8 njurbäckeninflammation
      4 njurbiopsi
      1 njurbipopsi
      6 njurcancer
      1 njurceller
      1 njurcellscarcinom
      1 njurdysfunktion
     10 njure
     26 njuren
      7 njurens
      1 njurepitelceller
      1 njurformade
      8 njurfunktion
      2 njurfunktionen
      1 njurglomeruli
      1 njurinfektion
      2 njurinflammation
      2 njurinsufficiens
      1 njurkomplikationer
      1 njurmissbildningar
      1 njurpåverkan
      2 njurproblem
      3 njursjuka
      7 njursjukdom
      3 njursjukdomar
      1 njursjukdoms
      1 njurskada
      7 njurskador
     14 njursten
      7 njurstenar
      1 njurstenenstenarna
     20 njursvikt
      1 njursvikten
      2 njursymtom
      3 njurtransplantation
      1 njurtransplantationen
      2 njurtubuli
      1 njurvävnaden
      5 njuta
      1 njuter
     12 njutning
      2 njutningen
      1 njutningskänsla
      4 njutningsmedel
      1 njutningsmedlen
      2 nkceller
      1 nkcellslymfom
      1 nkr
      1 nl
      1 nlm
      1 nlp
     11 nm
      1 nmda
      1 nmdaaktivitet
      1 nmdaantagonister
      3 nmdareceptorer
      1 nmdareceptorerna
      7 nmdareceptorn
      1 nmdareceptorns
      1 nmdareceptorstimulering
      1 nmdareceptorsubenheter
      1 nmdateorin
      2 nmoll
      1 nmranalyser
      1 nnrti
      1 �nns
     10 no
      1 noak
      1 nobel
      1 nobelförsamlingens
      8 nobelpris
      1 nobelprisbelönta
     19 nobelpriset
      2 nobelpristagare
      4 nobelpristagaren
      1 nobels
      1 nocardia
      2 nocebo
      1 noceboeffekt
      3 noceboeffekten
      1 nocere
      2 nociceptiv
      2 nociceptiva
      1 nociceptorerna
      1 nocturn
      1 nocturnus
      1 nöd
      1 nödår
      1 nödbromsning
      1 noddack
      1 noder
      2 nödfall
      1 nödig
      1 nödinsatser
      1 nödläge
      1 nödlösning
      3 nödnummer
      1 nödnumret
      3 nodosus
      1 nödrutschkana
      4 nödsituation
      1 nödsituationen
      4 nödsituationer
      1 nödslaktas
      1 nödsocker
      2 nödställda
      1 nödtillstånd
      2 nödtrakeotomi
      1 nödtvång
      1 noduliformation
      1 nödutgång
      3 nödutgångar
      1 nödutgången
      1 nödutrymning
     31 nödvändig
     16 nödvändiga
      1 nödvändiggöra
      1 nödvändighet
     48 nödvändigt
     32 nödvändigtvis
      2 noe
      2 noes
      1 noetiska
     23 nog
     11 noga
     19 noggrann
      7 noggranna
      3 noggrannare
      8 noggrannhet
      2 noggrannheten
     14 noggrant
      1 nogier
      1 nogsamt
      1 noirgenren
      1 noise
      3 nöja
      4 nöjda
      1 nöjde
      1 nöje
      1 nöjer
      1 nöjes
      2 nöjesdroger
      1 nöjesparker
      4 nokturi
      1 nokturn
      2 nolan
      7 noll
      1 nollresultat
      1 nollsummespel
      3 nollvision
      2 noma
      1 nomadiserade
      1 nomadiska
      2 nomenklatur
      1 nomenklaturen
      1 nominatunderarten
      1 nominell
      1 nominellt
      1 nominerades
      1 nominering
      1 nomos
      4 non
      1 nonapeptider
      1 noncaffeinated
      1 noncaloric
      1 nonchalant
      2 nonhodgkins
      1 nonie
      1 nonien
      2 noninvasiv
      1 nonsensord
      1 nonsuicidal
      5 nonylfenol
      1 nonylfenoletoxilater
      1 noomi
      1 noordbrabant
      1 nope
      1 nor
     18 noradrenalin
      2 noradrenalinet
      2 norberg
     12 nord
      2 nordafrika
     40 nordamerika
      3 nordamerikanska
      2 nordamerikas
      1 nordanvind
      1 nordanvinden
      2 nördar
     32 norden
      1 nordenfelt
      1 nordens
      5 nordeuropa
      1 nordeuropéernas
      1 nordeuropeisk
      1 nordhavsräka
      1 nördighet
     14 nordisk
     19 nordiska
      1 nordiske
      2 nordiskt
      1 norditalien
      1 nordlig
      3 nordligare
      1 nordligast
      2 nordligaste
      1 nordöstra
      1 nordsjön
      1 nordstedt
      1 nordström
      1 nordtyska
      1 nordvästeuropeisk
     12 nordvästra
      1 norell
      1 norepinefrin
     45 norge
      4 norges
      1 nori
      7 norm
    116 normal
    138 normala
      1 normalandel
      3 normalbefolkningen
      2 normalbegåvade
      3 normalbegåvning
      2 normalbelastad
      1 normalbyggda
      1 normalen
      1 normaler
      1 normalfall
      1 normalfallen
     13 normalfallet
      2 normalfärgad
     12 normalflora
      9 normalfloran
      1 normalflorans
      1 normalfördelad
      1 normalfördelade
      1 normalfördelning
      1 normalfördelningen
      1 normalfungerande
      1 normalfysiologin
      1 normalfysiologiska
      1 normalgräns
      1 normalgrupp
      1 normalhörande
      1 normalinställning
      1 normalisation
      2 normalisera
      1 normaliserad
      5 normaliseras
      1 normalisering
      1 normaliseringen
      7 normalitet
      1 normalläget
      2 normallång
      1 normallånga
      2 normallängd
      1 normallängden
      1 normalnivå
      1 normalpigmenterad
      2 normalpopulation
      7 normalpopulationen
      1 normalposition
      2 normalprocess
      1 normalpsykologi
      2 normalpsykologin
      1 normalspermiebildning
      1 normalställning
      2 normalstort
    346 normalt
      2 normaltillstånd
      1 normaltillståndet
      1 normaltryckshydrocefalus
      1 normalutveckling
      1 normalvärden
      2 normalvärdet
      2 normalvariationen
      1 normalvävnaden
      1 normalvikt
      3 normalviktig
      1 normalviktiga
      1 normalzonen
      4 norman
      1 normandisk
      1 normans
      2 normativa
      4 normen
     14 normer
      1 normera
      2 normerade
      1 normeringsgrupp
      1 normerna
      2 normgruppen
      2 normgruppens
      1 normlöshet
      3 normoblast
      1 normsystem
      1 norovirus
      1 noroviruset
      7 norr
     37 norra
      1 norrbotten
      1 norrbottens
      1 norrköping
      3 norrland
      4 norrlands
      1 norrlandsgränsen
      1 norrländsk
      1 norrländska
      1 norrländskt
      1 norrlandskusten
      1 norrmalmstorg
      1 norrmalmstorgsdramat
      2 norrmalmstorgssyndromet
      1 norrmän
      2 norrmannen
     10 norrut
      6 norsk
      6 norska
      1 norskan
      1 norskans
      2 norskt
      1 norsktfinskt
      3 north
      1 northern
      1 northwest
      1 norvasc
      1 norwalk
      1 norwalkinfektion
      3 nos
      1 nose
      1 nosen
      1 noskvalster
      1 nosokomiala
      6 nosologi
      2 nosologin
      1 nosomani
      1 nosos
      1 nosotras
      1 nosstyng
      6 not
      7 nöt
      5 nötallergi
      2 nötboskap
      3 noter
     13 notera
      3 noterade
      2 noterades
      1 noterar
     14 noteras
      3 noterat
      5 noterats
      1 noterbara
      2 noterbart
      2 noteringar
      1 nötfett
      1 nötfluga
      1 nötfria
      2 notis
      1 notiser
      1 nötkärnorna
     18 nötkreatur
      3 nötning
      1 notokord
      1 notoriska
      2 notoriskt
      1 nötrasen
      1 nötstyngen
      1 notte
     17 nötter
      7 nous
      5 nov
      1 nova
      1 novell
      1 noveller
     24 november
      1 novgorod
      1 novocain
      1 novokain
      1 novolizer
      1 novomedopa
      1 novopulmon
      1 novorapid
      1 novum
      2 np
      1 nph
     11 nr
      1 nrel
      1 nremsömn
      1 nrti
      2 nsa
     12 nsaid
      1 nsaider
      1 nsaidläkemedelsgruppen
      7 nsaidpreparat
      1 nsaids
      1 nsaidtyp
      1 nspot
     24 nssi
      3 nt
      2 nterminala
      1 nterminalen
      1 nterminalerna
      1 ntsc
    137 nu
      1 nubafolket
      1 nuc
      1 nuclear
      1 nucleus
      1 nudlar
      1 nuet
      1 nufers
      1 nuffield
      8 nuförtiden
      1 nugget
      1 nukleär
      2 nukleära
      2 nuklearmedicin
      1 nukleärmedicin
      1 nuklearmedicinsk
      2 nukleärmedicinsk
      1 nukleärmedicinska
      2 nukleinsyra
      2 nukleinsyraamplifiering
      1 nukleinsyradetektion
      1 nukleinsyradetektionstesterna
      1 nukleinsyrasyntes
      1 nukleinsyratest
      1 nukleinsyror
      1 nukleinsyrornas
      2 nukleofil
      1 nukleofila
      1 nukleofiler
      1 nukleokapsid
      1 nukleoler
      1 nukleosidanaloger
      1 nukleosider
      2 nukleotid
      1 nukleotider
      1 nukleotidsekvenser
      1 nukleotidsyntesen
      5 nuläget
      2 numer
    132 numera
      1 numeriska
      1 numeriskt
     12 nummer
      2 nummerkonto
      5 nummerkonton
      1 numrerade
      1 numreras
      1 numret
      1 nunna
      1 nunneörts
      1 nunnor
      2 nürnberg
      1 nürnbergkonventionen
      1 nürnbergrättegångarna
      2 nurse
      1 nursepatient
      3 nursing
      1 nursingtekniker
      1 nuss
      1 nussbaum
      4 nussmetoden
      1 nussoperationer
      9 nutida
     11 nutrition
      3 nutritionist
      1 nutritionisten
      2 nutritionistens
      3 nutritionister
      1 nutritionsforskningen
      1 nutritionskommitté
      1 nutritionslära
      2 nutritionsområdet
      1 nutritionsrubbningar
      1 nutritionsstörningar
     28 nuvarande
      1 nuvaring
      1 nuvenia
      1 nuxvomica
      6 nv
    125 ny
    267 nya
      1 nyandlighet
      5 nyans
      7 nyanser
      2 nyanserade
      1 nyanserar
      1 nyansskiftande
      1 nyansskillnader
      1 nyår
      1 nyara
     24 nyare
      1 nyårsafton
      1 nyaste
      1 nyberg
      1 nybildad
      3 nybildade
      1 nybildandet
      2 nybildas
     12 nybildning
      1 nybildningen
      1 nyblidning
      1 nyblivet
      6 nyblivna
      2 nybörjare
      1 nybörjares
      1 nybro
      1 nybyggnationer
      1 nycanders
      2 nyckel
      2 nyckelbenet
      1 nyckelceller
      1 nyckelexperimentet
      1 nyckelhålsliknande
      1 nyckelhålspupill
      1 nyckelknippa
      1 nyckelmotiv
      1 nyckeln
      2 nyckelord
      1 nyckelretningar
      2 nyckelroll
      2 nyckeltal
      1 nycomed
      1 nydestillerat
      1 nydiagnostiserade
      2 nyfiken
      4 nyfikenhet
      2 nyfödd
     33 nyfödda
      1 nyföddas
      1 nyförlöstas
      4 nyfött
      1 nygaard
      1 nygårds
      1 nygrekiska
      1 nyha
      3 nyhet
      3 nyheter
      1 nyheterna
      1 nyhetsbrev
      1 nyhetskaraktär
      1 nyhetsprogram
      1 nyhetssändning
      1 nyinrättade
      1 nyinsatta
      3 nykläckta
      3 nykter
      1 nykterhet
      1 nyktra
      1 nyktrat
      1 nyktre
      1 nyktres
      2 nykturi
      1 nyland
      3 nylat
      5 nylatin
      2 nylatinets
      1 nylatinska
     40 nyligen
      6 nylon
      1 nylonmembran
      1 nylonteflon
      1 nymalthusianismen
      1 nymåne
      1 nymf
      1 nymfen
      4 nymfer
      2 nymutation
      1 nymutationer
      1 nyopererad
      2 nypa
      1 nyplatonismen
      1 nyps
      1 nyquistteoremet
      1 nyrekrytering
      1 nysa
      1 nyse
      4 nyser
      1 nyses
      1 nyskrivna
      7 nysning
      7 nysningar
      4 nysningen
      1 nysört
      1 nysrotsväxter
      3 nyss
      1 nyssnämnda
      6 nystagmus
      1 nytänkande
      1 nytestamentliga
      1 nytillväxt
      1 nytryck
     45 nytt
     32 nytta
     11 nyttan
      1 nyttavsnittlÄnk
      5 nyttig
     12 nyttiga
      4 nyttigt
      3 nyttja
      1 nyttjad
      1 nyttjade
      1 nyttjades
      2 nyttjar
      2 nyttjas
      1 nytto
      4 nyttobakterier
      1 nyttobakterierna
      1 nyttodjur
      2 nytvättade
      1 nyupptäckt
      1 nyupptäckta
      1 nyutvecklad
      1 nyväckta
      1 nyvitalism
      1 nyvunnen
      2 nyzeeländske
      1 nzara
     17 o
      2 �ó
      1 ���ó
      1 ����ó
      4 ö
      1 Ö
      1 oacceptabelt
      3 oacceptabla
      1 oaccepterad
      2 oaccepterat
      1 oädel
      1 oae
      3 oak
      1 oakdermatit
      1 oakley
      2 oäkta
      1 oaktat
      1 oändlig
      1 oändligt
      2 oangenäm
      2 oansenligt
      1 oansvarigt
      1 oanvänd
      1 oanvändbar
      2 oanvändbara
      9 öar
      7 öarna
      1 oartig
      1 oas
      1 oaspirerad
      2 oaspirerade
      2 oaspirerat
      1 oat
      1 oåterkallelig
      1 oåterkalleliga
      1 oåterkalleligt
      1 oates
      2 oätlig
      1 oattraktivt
      3 oavbrutet
      1 oavbrutna
      1 oavhängigt
     44 oavsett
      1 oavsiktlig
      3 oavsiktligt
     22 obalans
      1 obalansen
      1 obalanser
      1 obalanserad
      1 obalanserat
      1 obducerade
      1 obducerat
      1 obducerats
      1 obduco
      1 obductio
     10 obduktion
      7 obduktioner
      1 obduktionsfynd
      1 obduktionssalarna
      4 obefintlig
      3 obefintliga
      3 obefogad
      1 obefogat
      3 obefruktade
      1 obefruktat
      1 obegränsad
      1 obegripligt
     34 obehag
      2 obehagen
      1 obehaget
     14 obehaglig
     16 obehagliga
     12 obehagligt
      2 obehagskänslor
      1 obehagsproducerande
      1 obehagströskel
      2 obehagströskeln
     40 obehandlad
     13 obehandlade
     16 obehandlat
      1 obehindrat
      1 obehörig
      1 obehöriga
      1 obehörigen
      2 obekräftade
      3 obekväm
      4 obekväma
      3 obekvämt
      1 obekymrat
      1 obemannad
      2 obemärkt
      1 obemärkta
      1 obenägna
      1 obenthet
      1 obeprövade
      1 oberfruktade
     51 oberoende
      1 oberörda
      1 obesatta
      1 obesefetma
      1 obesitas
      1 obesity
      1 obesläktad
      1 obesvärad
      1 obesvärat
      2 obetalda
      1 obetingat
      1 obetvinglig
      2 obetvingliga
      1 obetvingligt
      3 obetydlig
      1 obetydliga
      3 obetydligt
      1 obevakade
      1 obevekligt
      1 obevisade
      1 obevisat
      1 obildad
      1 obildbara
      1 object
     50 objekt
     25 objektet
      5 objektiv
      6 objektiva
      1 objektivism
      9 objektivt
      1 objektrelation
      2 objektrelationer
      1 objektrelationsskolan
      3 objektrelationsteori
      5 objektrelationsteorin
      1 objektrelationsteorins
      2 oblekt
      1 oblektofärgat
      1 obligata
      4 obligationer
      1 obligationerna
      2 obligatorisk
      1 obligatoriska
      6 obligatoriskt
      2 obliquus
      1 obliterans
      5 oblongata
      1 oboens
      3 obotlig
      2 obotligt
      1 obrännbart
      1 obrien
      1 obrukbar
      2 obrukbart
      2 obrutna
      1 obscena
      1 obscent
      1 observans
      1 observant
      9 observation
      1 observational
     15 observationer
      1 observationsförmåga
      1 observationskategorier
      1 observationsmaterial
      1 observationstuben
      1 observatör
      1 observatörsstatus
     18 observera
      7 observerade
      2 observerades
      4 observerar
     15 observeras
     12 observerat
      7 observerats
      1 observerbar
      1 observerbara
      1 obsessioner
      1 obsessive
      1 obsessivecompulsive
      2 obsidian
      1 obsolet
      1 obsoleta
      1 obstetricia
      4 obstetrik
      1 obstetriken
      1 obstetrikens
      2 obstetriker
      1 obstetrisk
      1 obstetriska
      2 obstetrix
      1 obstipation
     10 obstruktion
      1 obstruktionen
     15 obstruktiv
      6 obstruktiva
      1 obstruktivt
      1 obtusata
      1 oc
      2 ocampa
      1 ocampierna
      1 occh
      1 occidentalis
      1 occipational
      1 occludiner
      1 occulta
      1 occupation
     11 occupational
      1 occurrence
     16 ocd
      3 ocdpatienter
      1 ocdsymptom
      1 oceanografi
  21749 och
      1 ochangiodysplasi
      1 ochblododlingar
     93 ocheller
      1 ochlerotatus
      1 ochmaskar
      1 ochökad
      1 ochroleucus
      1 ochrus
      1 ockelbo
      3 ockelbosjuka
      3 ockelbosjukan
      1 ockelboviruset
      1 ockham
      1 ockluderingsanordning
      1 ocklusion
      1 ockra
   1659 också
      1 ockult
      1 ockupationen
      1 ockuperas
      1 ocn
      2 oconnor
      1 octavianus
      1 ocular
      1 ocularist
      1 ocularists
      1 oculomotoriuspares
      5 odd
      1 oddi
      3 oddskvot
      2 oddskvoten
      1 oddskvoterna
      1 oddskvoternas
      5 öde
      1 ödegårdsprojektet
      1 ödeläggande
      2 odelbar
      1 odelbara
     23 ödem
      4 Ödem
      1 ödembildning
      1 ödemen
      1 Ödemet
      2 oden
      1 odense
      1 odenwald
      2 ödesdigert
      2 ödesdigra
      1 ödesgudinnorna
      1 ödets
      1 odiagnostiserat
      5 odifferentierad
      1 odifferentierade
      1 odiskutabelt
      1 odjuret
     12 odla
      3 ödla
      3 odlad
     15 odlade
      3 odlades
      3 ödlan
      2 ödlans
     35 odlas
      4 odlats
      1 ödlefamiljen
      1 ödlekött
      3 ödleungarna
     19 odling
      2 odlingar
      1 odlingsbehållaren
      1 odlingsdiagnostik
      1 odlingsformen
      1 odlingskulturens
      1 odlingsområdena
      1 odlingsprov
      1 odlingstest
      1 odlingszon
      6 ödlor
      1 ödlorna
      1 ödlornas
      1 Ödlornas
      1 ödmjuka
      5 odödlighet
      1 odödligheten
      2 odone
      1 odontofobi
      3 odontologi
      3 odontologie
      2 odontologin
      8 odontologisk
      4 odontologiska
      4 odör
      1 odp
      1 odrickbar
      1 odugliga
      1 odysseus
      1 oecdländerna
      1 oecdnea
      1 oecds
      1 oedema
      1 oeftergivlig
      1 oeftergivliga
      1 oeftergivligt
      5 oegentligt
      1 œillet
      1 oelastisk
      1 oemotståndlig
      1 oengagerad
      1 oengagerat
      4 oenighet
      1 oenigheter
      2 oerfarna
      8 oerhört
      1 oersättliga
      1 oesophagus
      2 oestetiska
      1 oestridae
      1 oestring
      1 oestrus
    148 of
      1 ofäränderlig
      1 ofärgat
     22 ofarlig
     22 ofarliga
      1 ofarlighet
     16 ofarligt
      1 ofarrell
      2 ofelbart
      1 offensiv
      1 offensiva
      1 offensiven
      1 offensivt
     15 offentlig
     39 offentliga
      1 offentligas
      1 offentliggjorde
      1 offentlighetsprincipen
      9 offentligt
     31 offer
      1 offerhåvarna
      1 offertoriet
      1 offerviljan
      1 office
      1 officerare
      8 officiell
     10 officiella
     18 officiellt
      4 officinalis
      1 officinarum
      1 offrades
      1 offrar
      1 offrats
      9 offren
      1 offrens
     11 offret
      3 offrets
      1 ofint
      1 ofixerat
      4 ofödda
      1 oföränderlig
      1 oföränderliga
      2 oföränderligt
      1 oförändlighet
      8 oförändrad
      3 oförändrade
      5 oförändrat
      1 oförargliga
      1 oförargligt
      1 oförberett
      1 oförbrända
      2 ofördelaktig
      2 oförenliga
      1 oförklarat
      1 oförklarlig
      1 oförklarliga
      3 oförklarligt
      1 oförlösta
     40 oförmåga
      1 oförmågaallergi
      2 oförmågan
      7 oförmögen
      1 oförmöget
      1 oförmögna
      1 oförskriven
      1 oförståeliga
      1 oförståelse
      1 oförstörande
      1 oförstörlbar
      1 oförtjänt
      2 oförutsägbar
      3 oförutsägbara
      2 oförutsägbart
      2 oförutsedda
      1 ofött
      1 ofrånkomliga
      1 ofri
     10 ofrivillig
     14 ofrivilliga
     11 ofrivilligt
      1 ofruktsamhet
   1543 ofta
      2 oftalmiska
      1 oftalmolog
      1 oftalmologassistenter
      1 oftalmologer
      2 oftalmologi
      1 oftalmologin
      1 oftalmologiska
      1 oftalmomyiasis
      6 oftalmoskop
      2 oftalmoskopet
     67 oftare
    631 oftast
      1 oftats
     12 ofullständig
      1 ofullständiga
      1 ofullständigt
      1 ofullvärdiga
      1 öfvade
     25 öga
      1 ögas
      2 ogästvänlig
      1 ogästvänliga
     79 ögat
      1 ögathjärnan
     29 ögats
      1 Ögats
      2 ogenomtränglighet
      2 ogenomträngligt
      4 ogift
      7 ogifta
      3 ogifte
      1 ogiftig
      3 ogiftiga
      3 ogillar
      2 ogiltigt
     44 ögon
      2 ögonbindel
      2 Ögonbindel
      3 ögonblick
      1 ögonblickets
      1 ögonblickliga
      1 ögonblickligen
      3 ögonbotten
      5 ögonbryn
      2 ögonbrynen
      1 ögonbrynsbåge
      1 ögonbrynsben
      1 ögondarrning
      2 ögondiagnostik
      1 Ögondiagnostik
      5 ögondroppar
      2 Ögondroppar
      1 ögoneffekten
     72 ögonen
      2 Ögonen
      4 ögonens
      4 ögonfärg
      1 ögonfärgen
      3 ögonfransar
      5 ögonfransarna
      1 ögonglob
      2 ögongloben
      1 ögonglober
      1 ögonhåla
      2 ögonhålan
      1 ögonhålen
      2 ögoninfektion
      1 ögonirritation
      2 ögonkirurgi
      1 ögonklotet
      2 ögonkontakt
      1 Ögonkontakt
      9 ögonläkare
      1 ögonläkaren
      1 ögonlapp
      1 Ögonlappar
      1 ögonlaserkirurgin
      1 ögonlins
      8 ögonlock
      5 ögonlocken
      8 ögonlocket
      1 ögonlockets
      1 ögonlockshygien
      1 ögonlocksinflammation
      1 ögonlockskanterna
      1 ögonmissbildning
      1 ögonmuskelstörningar
      1 ögonmusklerna
      1 ögononkologiska
      2 ögonöppning
      1 Ögonöppning
      1 ögonoptik
      1 ögonpatologiska
      4 ögonproblem
      2 ögonprotes
      4 ögonproteser
      1 Ögonproteser
      1 Ögonproteserna
      1 ögonreaktioner
      1 ögonregionen
      1 ögonretande
     12 ögonrörelser
      3 ögonrörelserna
      1 ögonrörelserubbningar
      1 ögonrörlighet
      3 ögonsjukdom
      4 ögonsjukdomar
      3 Ögonsjukdomar
      2 ögonsjukdomen
      1 ögonsjuksköterskor
      1 ögonskada
      2 ögonskador
      1 ögonskugga
      1 Ögonskugga
      1 ögonskuggor
      1 Ögonskuggor
      1 Ögonspegel
      2 ögontryck
      1 Ögontryck
      1 ögonundersökning
      4 ögonvitor
      2 ögonvitorna
      1 Ögonvitorna
      1 ögonvrån
      6 ogräs
      1 ogräsfrön
      2 ogräsmedel
      1 ogrenad
      3 ogrenade
      4 ogynnsam
      6 ogynnsamma
      3 ogynnsamt
      3 oh
      1 ohållbar
     43 ohälsa
      1 ohälsan
      3 ohälsosam
      1 ohälsosamma
      1 ohälsotillstånd
      2 ohämmad
      1 ohämmat
      1 ohanterlig
      1 ohara
      1 ohbindande
      1 ohda
      2 ohgrupp
      5 ohgruppen
      2 ohgrupper
      2 ohgrupperna
      2 ohio
      1 Öhman
      1 ohmmeter
      1 ohmolekylen
      1 ohms
      2 ohne
      1 ohövlig
      1 ohsas
      1 ohydrerade
      1 ohyfsat
      1 oidentifierad
      1 oidentifierade
      1 oidipus
      2 oidipusmyten
      1 oigenkännlighet
      1 oinfekterade
      1 oinsatte
      1 ointelligent
      1 ointelligenta
      2 ointressant
      1 ointressanta
      1 ointresserad
      1 ojämförligt
      1 ojämlikhet
      4 ojämn
      1 ojämna
      1 ojämnare
      2 ojämnhet
      5 ojämnheter
      1 ojämnt
      1 ok
    138 öka
    205 ökad
      9 Ökad
     87 ökade
      2 Ökade
     34 okänd
      1 ökänd
     13 okända
      2 ökända
      1 okändas
     22 ökande
      1 Ökandet
      1 okändref
      1 okänslig
      1 okänsliga
      2 okänslighet
     17 okänt
    339 ökar
      9 ökas
    110 ökat
      5 Ökat
      1 okay
      1 okej
      1 ökenödla
      2 ökenområden
      1 ökentaipan
      1 oklädda
      1 oklahoma
      1 oklanderligt
     13 oklar
      5 oklara
      2 oklarheter
     32 oklart
      1 oklassificerbara
      1 oklorfenol
      3 öknamn
      1 öknamnet
      1 okning
     51 ökning
      1 Ökning
      1 ökningar
     19 ökningen
      5 Ökningen
      2 okokt
      5 okomplicerad
      3 okomplicerade
      1 okomplicerat
      1 okoncentrerad
      1 okoncentrerat
      9 okontrollerad
      1 okontrollerade
      9 okontrollerat
      3 okontrollerbar
      1 okontrollerbara
      1 okontrollerbart
      1 okontroversiellt
      1 okonventionella
      1 okorrigerad
      1 okritisk
      1 okritiskt
      1 oktan
      1 oktantal
      4 oktav
      1 oktettregeln
     21 oktober
      1 oktoberstormhatt
      1 okular
      1 okulär
      1 okulära
      1 okularist
      2 okularister
      1 okunnig
      1 okunnighet
      3 okunskap
      1 okvalificerade
      1 ol
      8 öl
      1 oladdade
      1 olag
      2 olaga
      1 olägenhet
      1 olägenheter
      2 olaglig
      3 olagliga
     14 olagligt
      5 olämplig
      5 olämpliga
      9 olämpligt
      7 Öland
      1 olanzapin
      1 oläsbara
      2 ölbryggning
      1 old
      1 ole
      9 oleander
      4 oleanderväxter
      1 oledade
      1 olekranonbursit
      1 olevande
      1 olfactorius
      1 olfaktorisk
      1 olfaktoriska
      1 oligofruktos
      1 oligomer
      2 oligonukleotid
      1 oligosackarider
      1 oligozoospermi
      4 oliguri
      5 olik
   1699 olika
      3 olikartade
      2 olikartat
      1 olikfärgade
      1 olikhet
      6 olikheter
      1 olikheterna
      1 olikpoliga
      3 olikt
      2 olivecrona
      1 olivecronas
      1 oliver
      1 olivgrön
      1 olivgrönt
      1 olivier
      5 olivolja
     22 olja
      8 oljan
      1 oljans
      1 oljebaserade
      1 oljebaserat
      1 oljefärger
      1 oljeinnehåll
      1 oljekanaler
      1 oljekylning
      1 oljepalmen
      1 oljesyra
      1 öljett
      1 öljetten
      1 öljetter
      1 Öljetter
      1 oljeväxter
      2 oljig
      1 oljiga
     19 oljor
      7 oljorna
      1 oljornas
      4 oljud
      1 oljudet
      3 olle
     19 ollonet
      1 ollonkanten
      4 olof
      1 olofsson
      1 ologiska
      2 ologiskt
      1 olönsamt
      4 olöslig
      9 olösliga
      8 olösligt
      1 olöst
      2 olovlig
      4 olsson
      2 olust
     14 olycka
      8 olyckan
      2 olycklig
      4 olyckliga
      1 olyckligt
     26 olyckor
      3 olyckorna
      1 olycks
      1 olycksdiger
      9 olycksfall
      1 olycksfallen
      3 olyckshändelse
      1 olycksorsaker
      2 olycksplats
      1 olycksrelaterade
      1 olycksrisker
      3 olympiska
      1 olympiske
   3299 om
      9 öm
      2 oma
      2 omalizumab
      1 omanlig
      1 omanliga
      1 omarbetats
      1 omärkt
      1 omasum
      1 omätbar
      3 omätbara
      1 omättade
      1 omättat
      1 omättnaden
      1 ombads
      1 ombesörjs
      1 ombetäckningar
      1 ombilda
      1 ombildad
      5 ombildade
      1 ombildades
      3 ombildar
      7 ombildas
      1 ombildats
      5 ombord
      1 ombud
      1 ombyggnad
      1 ombyggnaden
      1 ombyggnadstiden
      1 omdebatterad
      1 omdebatterade
      2 omdebatterat
      1 omdirigeras
      2 omdiskuterad
      3 omdiskuterade
      1 omdiskuteras
      8 omdiskuterat
      5 omdöme
      1 omdömen
     29 omedelbar
      3 omedelbara
     30 omedelbart
      9 omedveten
      1 omedvetenhet
      8 omedvetet
     24 omedvetna
      1 omedvetnas
      9 omega
      1 omegafett
      1 omegafetter
      3 omegafettsyror
      1 omegafettsyrors
      1 omegafettysyror
      2 omeprazol
      1 ometyl
      1 ometylensubstituerade
      1 omfamnat
      2 omfång
      1 omfångsrika
     10 omfatta
     10 omfattade
     94 omfattande
     92 omfattar
     15 omfattas
      3 omfattat
     30 omfattning
      4 omfattningen
      1 omflyttning
      1 omföderskor
      1 omfördelas
      1 omforma
      1 omformade
      1 omformas
      1 omformats
      1 omformulerat
      5 omgående
      4 omgång
      6 omgångar
      1 omgärdad
      1 omgärdar
      1 omgav
     18 omger
      5 omges
     50 omgivande
      2 omgiven
      3 omgivet
      4 omgivna
      1 omgivnade
     33 omgivning
      2 omgivningarna
     66 omgivningen
      1 omgivningenbr
      4 omgivningens
      4 omgivningsljud
      1 omgivningsradiologi
      1 omgivningstemperaturen
      1 omgivningstrycket
      1 omhänderta
     12 omhändertagande
      3 omhändertagandet
      1 omhändertas
     10 ömhet
      1 ömheten
      1 ömhetsbetygelser
      1 omhuldades
      1 omhuldat
      1 omkastning
      5 omkom
      1 omkommer
      2 omkommit
      1 omkomna
      1 omkopplingen
      3 omkrets
      2 omkretsen
    245 omkring
      6 omkringliggande
      2 omkringvarande
      1 omkullkastar
      1 omlades
      1 omlagda
      1 omläggningar
      1 omläggningen
      1 omlagras
      2 omlöpningar
      5 omlopp
      5 ömma
      1 ommålning
      7 ömmande
      1 ömmar
      1 ommayabehållare
      1 ommikroorganismer
      2 omnämnande
      1 omnämnanden
      4 omnämnd
      1 omnämnda
      2 omnämner
     12 omnämns
      1 omnär
      1 omnejd
      1 omnipotenta
      1 omniscienta
      1 omodernt
      1 omogen
      8 omogna
      4 omöjlig
      3 omöjliga
      1 omöjliggöra
      3 omöjliggörs
     24 omöjligt
      1 omoral
      3 omoraliskt
      1 omorganisation
      2 omorganiserades
      1 omorganiserar
      1 omorientering
      1 omotiverad
      1 omotiverade
      1 omött
      1 omöversatt
      1 omplacering
      1 omprioritering
      1 omprövat
      1 omprövningar
     93 område
    184 områden
     23 områdena
      1 områdenas
    119 området
      2 områdets
      1 omräknar
      1 omreglera
      1 omringar
      1 omritning
      3 omritningen
      2 omröstning
      1 ömsa
      1 ömsade
      1 omsänder
      2 ömsar
      1 omsätta
      1 omsättas
      2 omsätter
      4 omsättning
      8 omsättningen
      1 omsättningsbara
      2 omsätts
      4 ömsesidig
      1 ömsesidiga
      6 ömsesidigt
      1 omskakande
      1 omskakning
      2 omskärelse
      1 omskärning
      1 omskhemorragiskt
      1 omskriven
      1 omskrivet
      1 omskrivna
      2 omskrivning
      1 omskuren
      2 omskurna
      1 omslag
      1 omslutande
      5 omsluter
      1 omslutna
      2 ömsom
     18 omsorg
      1 omsorgen
      1 omsorger
      1 omsorgsarbete
      1 omsorgsförmåga
      3 omsorgsfullt
      1 omsorgslagen
      1 omsorgspersonalen
      1 omsorgspersoner
      2 omsorgsprogrammet
      1 omsorgsrationalitet
      3 omsorgstagare
      2 omsorgstagarna
      1 omsorgsvården
      1 omsorgsverksamheter
      1 omställning
     27 omständigheter
      3 omständigheterna
      1 omständlig
      1 omständliga
      1 omstörtande
      3 omstridd
      1 omstridda
      1 omstritt
      1 omstrukturerar
      1 omstruktureringen
      2 omsvängning
      4 ömt
      2 omtalade
      4 omtalas
      3 omtalat
      1 ömtålig
      2 ömtåliga
      1 omtanke
      1 omtöcknad
      3 omtöcknat
      1 omtolkade
      5 omtvistad
      1 omtvistade
      2 omtvistat
      5 omtyckt
      1 omtyckta
      1 omvägen
      2 omvälvande
      7 omvänd
      1 omvända
      1 omvändelse
     11 omvandla
      1 omvandlade
      1 omvandlades
     11 omvandlar
     51 omvandlas
      1 omvandlat
      2 omvandlats
      7 omvandling
      1 omvandlingar
      8 omvandlingen
      1 omvandlingsprodukt
      1 omvandlingstiden
      6 omvänt
      1 omvårdande
      3 omvärderande
      1 omvärdering
     13 omvårdnad
      4 omvårdnaden
      2 omvårdnadsdokumentation
      2 omvårdnadsforskning
      1 omvårdnadsforskningen
      1 omvårdnadspersoner
      1 omvårdnadsprofesstionen
      1 omvårdnadsprogrammet
      1 omvårdnadssocial
      1 omvårdnadssystem
      1 omvårdnadssystemet
      1 omvårdnadsteori
      1 omvårdnadsteorier
      1 omvårdnanden
      3 omvärld
     12 omvärlden
      2 omvärldens
      1 omvärldskunskap
      2 omväxlande
      2 omyndig
      3 omyndiga
      1 omyndigförklara
     25 on
      4 ön
      1 onan
      1 onanerar
      1 onani
      1 önationer
      2 onaturlig
      2 onaturliga
      4 onaturligt
      1 onchocerca
      2 onchocerciasis
      5 ond
     14 onda
      1 onde
      1 ondes
      1 ondines
      1 ondska
      1 ondskan
      1 one
      1 Önh
      1 Önhklinik
      2 onkgener
      5 onkogen
      2 onkogena
      6 onkogener
      4 onkologi
      2 onkologiska
      1 ónkos
      1 onliehtan
      3 online
      1 onlineaffärer
      1 only
      1 ono
      4 onödan
      5 onödig
      1 onödiga
      6 onödigt
     18 onormal
     13 onormala
     26 onormalt
      1 onormaltelektrokardiogram
      1 onsdagen
      1 onsenal
      2 onset
      3 önska
      3 önskad
     12 önskade
      6 önskan
     20 önskar
      1 Önskar
      3 önskas
      6 önskat
      4 önskemål
      2 önskningar
      5 önskvärd
      6 önskvärda
     10 önskvärt
     52 ont
      1 ontologisk
      1 ontologiska
      1 oocysta
      1 oocystor
      1 oocystorna
      1 oocyt
      1 oocyten
      2 oocyter
      1 oogama
      1 oogami
      1 oogenes
      1 oogenesen
      2 ookinet
      1 oomskurna
      1 oomyceten
      7 oönskad
     14 oönskade
      5 oönskat
      1 oönskvärda
      1 oöppnad
      2 oordnat
      2 oordning
      2 oorganisk
      3 oorganiska
      1 oorganiskt
      1 oosporer
      1 �o�ox
      1 ooxiderat
      1 op
      1 opaciteter
      2 opal
      2 opålitlig
      1 opålitliga
      1 opaproteinerna
      1 oparfymerad
      1 oparfyrmerat
      1 oparig
      3 opassande
      1 opastöriserad
      1 opastöriserade
      2 opåverkad
      2 opåverkade
      1 opera
      6 operant
      1 operarad
    121 operation
     58 operationen
      1 operationens
     49 operationer
      2 operationerna
      1 operationernas
      1 operationsärret
      2 operationsavdelning
      1 operationsavdelningen
      1 operationsbord
      1 operationsgruppen
      1 operationshålet
      1 operationsläran
      3 operationsmetod
      2 operationsmetoden
      2 operationsområdet
      1 operationsresultatet
      1 operationsresurser
      1 operationssalar
      1 operationssalarna
      1 operationssnitt
      1 operationsteknik
      1 operationstekniken
      2 operativ
      6 operativa
      1 operativsystem
      3 operativt
      1 opératoire
      1 operatören
      1 operatörens
     18 operera
      1 opererad
      7 opererade
      3 opererades
      1 opererande
     11 opererar
     30 opereras
      2 opererat
      2 opererats
      1 operforerat
      1 opersonliga
      1 ophiophagus
      1 ophthalmos
      1 opi
      2 opiat
      1 opiatberoende
      9 opiater
      1 opiatmissbruk
      1 opiatmissbrukare
      1 opiatmissbrukaren
      1 opigmenterade
      1 opii
      1 opinion
      1 opinionsbildningmalaria
      1 opinionsundersökningsföretaget
      1 opioiden
     12 opioider
      1 opioidpreparatmorfinderivat
      1 opioidreceptorer
      1 opioidsystemet
      1 opiopeptid
     11 opium
      1 opiumdroppar
      2 opiumhålorna
      1 opiumkrigen
      1 opiumrökandet
      2 opiumrökning
      3 oplanerade
      1 oplanerat
      1 opolär
      1 opolära
      1 opolärt
     23 öppen
      2 Öppen
      1 öppenhet
      1 öppenheten
     10 öppenvård
      1 Öppenvård
      6 öppenvården
      1 öppenvårdsapotek
      1 öppenvårdsbehandling
      2 öppenvårdsenheter
      1 öppenvinkelglaukom
     14 öppet
      1 öppetstående
     34 öppna
      1 Öppna
      1 öppnad
     14 öppnade
      2 Öppnade
      7 öppnades
      1 Öppnande
      1 öppnandet
     14 öppnar
     25 öppnas
      3 öppnat
      4 öppnats
     22 öppning
      4 öppningar
      1 öppningarna
      6 öppningen
      1 Öppningen
      1 öppningmun
      2 öppningsbar
      1 öppningsbara
      1 öppningsceremonin
      3 öppningsgrad
      1 öppningstid
      1 öppningstrycket
      1 opponerade
      1 opportunism
      2 opportunister
      4 opportunistiska
      1 opposites
      2 opposition
      1 oppositional
      1 oppositionen
      1 opraktiskt
      2 oprecis
      1 opressade
      2 oproblematiskt
      1 oproportionella
      1 oproportionerligt
      2 oprövade
      1 oprovocerade
      1 opsis
      1 opsonisering
      3 optik
     16 optiker
      1 optikerförbundet
      1 optikerförbundets
      5 optikern
      2 optikerna
      1 optikeroptometrist
      1 optikers
      1 optikuskolobom
      7 optimal
      7 optimala
     10 optimalt
      2 optimera
      2 optimering
     14 optimism
      1 optimismbias
      1 optimismen
      1 optimisten
      3 optimister
      1 optimistiska
      1 option
      3 optisk
     13 optiska
      8 optiskt
      1 optometri
      1 optotyper
      2 optotyperna
      1 optyl
      1 opubicerade
      4 or
      1 �ór
      1 ora
      8 öra
      1 oraffinerade
      1 oraffinerat
      1 orahilly
      1 oraklet
     28 oral
     14 orala
      1 oralazitromycin
      1 oralkirurgi
      1 oralmotorisk
      7 oralsex
     10 oralt
      8 orange
      1 orangegula
      1 orangeröda
      1 orangutanger
     30 örat
      2 oratium
      6 örats
      1 orätt
      2 orättvis
      2 orättvisa
      3 orättvist
      1 orbitan
      1 orbitofrontalcortex
      3 orcenia
      1 orchidopexi
      1 orchis
    110 ord
      1 ordagranna
      7 ordagrant
      1 ordavkodning
      2 ordavkodningen
      1 ordbehandla
      1 ordbilder
      1 ordblindhet
      1 ordböcker
      1 ordbok
      1 orddelar
     23 orden
      1 ordens
      6 ordentlig
      1 ordentliga
     24 ordentligt
      6 order
    227 ordet
      5 ordets
      4 ordförande
      1 ordförråd
      1 ordförrådet
      1 ordförrådsbaserade
      1 ordglömska
      1 ordinära
      5 ordinarie
      4 ordination
      2 ordinationen
      3 ordinera
      2 ordinerad
      1 ordinerade
      5 ordinerar
     19 ordineras
      1 ordinerat
      1 ordines
      1 ordkombination
      1 ördmedicin
      4 ordna
      1 ordnad
      6 ordnade
      1 ordnar
      2 ordnas
      1 ordnat
     31 ordning
      1 ordningar
     22 ordningen
      1 ordningsföljd
      1 ordningslagen
      1 ordningsproblem
      3 ordningsvakter
      2 ords
      2 ordsallad
      1 ordspel
      1 ordspråk
      1 ordstammen
      1 öre
      3 orealistiska
      8 Örebro
      8 oregelbunden
      1 oregelbundenhet
      1 oregelbundet
      8 oregelbundna
      1 oregerligt
      1 oreglerad
      1 oreglerat
      1 orelaterad
      1 orelaterat
      1 oren
      2 orena
      1 orenade
      1 orenat
      1 orencia
      2 orenheter
      1 orent
      1 oreserverade
      6 oresorberbara
      1 oresponsiv
     12 orexin
      1 orexinet
      1 orexininnehållande
      1 orexinliknande
      2 orexinnivåerna
      1 orexinreceptorer
      1 orfiril
    215 organ
      1 organbildningen
      2 organdonationer
      1 organdonatorn
      1 organdysfunktion
      1 organell
      3 organeller
     21 organen
      2 organens
     15 organet
      2 organets
      1 organett
      1 organförsämring
      2 organförstoring
      1 organfunktionen
      1 organhandel
      1 organicum
     32 organisation
     15 organisationen
      3 organisationens
     23 organisationer
      1 organisationerna
      1 organisationernas
      1 organisationers
      2 organisations
      2 organisationsförmåga
      1 organisationskonsulter
      1 organisationsmodellen
      2 organisationspsykologi
      2 organisationsutveckling
      3 organisatoriska
      4 organisera
      3 organiserad
      7 organiserade
      1 organiserande
      7 organiserar
      7 organiseras
      1 organiserat
      1 organisering
      1 organiseringen
     47 organisk
     58 organiska
     20 organiskt
     31 organism
     19 organismen
      7 organismens
     69 organismer
      7 organismerna
      3 organismers
      3 organisms
      3 organization
      1 organnivå
      1 organofosfat
      1 organogenesen
      6 organomegali
      1 organskador
      1 organstruktur
      3 organsvikt
     13 organsystem
      1 organsystemet
      3 organtransplantation
      1 organtransplantationer
      1 organviktsfaktorer
      1 organviktsfaktorn
     12 orgasm
      1 orgasmen
      1 orgasmens
      1 orgasmnjutning
      1 orgasmstörning
      1 orgastiska
      1 Örhänge
      7 örhängen
      2 Örhängen
      1 örhängesplaceringar
      1 örhänget
      1 Örhänget
      1 Örhängets
      1 orientalisk
      1 orientalism
      1 orientens
      5 orientera
      6 orienterad
      2 orienterade
      1 orienterat
      3 orientering
      1 orienteringstavlor
      1 origin
      3 original
      3 originalet
      1 originalmanus
      2 originalobservationer
      1 originalstudier
      2 originaltitel
      1 oriktiga
      3 oriktigt
      3 orimlig
      4 orimligt
      1 oripavin
      1 oripiment
      1 oris
      2 ork
      3 orka
      1 orkaner
     11 orkar
      2 orken
      1 orkeslös
      7 orkeslöshet
      1 orkestermedlemmarna
      1 orkestermusiker
      1 orkidéerna
      1 orksakar
      2 örlogsfartyg
      1 örlogsman
      8 orm
      1 orma
     18 ormar
      1 ormarna
      1 ormars
      1 ormartens
      1 ormarter
      1 ormarters
      1 ormattribut
      3 ormbär
      1 ormbärsörten
      7 ormbett
      1 ormbunkar
      3 ormbunksväxter
      9 ormen
      5 ormens
      1 ormfobi
      1 ormfobiker
      2 ormgestalt
      5 ormgift
      4 ormgifter
      1 ormgifters
      1 ormgiftsproducerande
      1 ormgudinnan
      1 ormkött
      1 ormlikt
      1 ormrotsflockelssläktet
      1 ormskinn
      1 ormvärlden
      2 ornament
      2 ornamenterade
      1 ornerade
      1 Örnhagen
      2 ornish
      1 ornithos
     48 oro
      2 oroa
      1 oroande
      1 orobus
      1 orofacial
      1 orofarynx
      7 orolig
      4 oroliga
      1 orolighet
      1 oroligt
      8 oron
     19 öron
      3 öronakupunktur
      2 öronbarn
      1 örondroppar
     27 öronen
      1 öronformad
      1 örongången
      1 öronhål
      1 öroninfektion
      2 öroninfektioner
     11 öroninflammation
      3 Öroninflammation
      4 öroninflammationer
      1 öroninsats
      2 öronkanalen
      1 öronkurett
      1 öronläkare
      9 öronljus
      2 Öronljus
      2 öronmusslan
      2 öronnäsahals
      1 öronnäsahalsläkare
      1 öronnäsahalssjukdomar
      2 öronproppar
      1 öronproteser
      1 öronsjukdom
      2 öronskabb
      2 Öronskabb
      1 öronskador
      2 öronsmärta
      2 öronsnäckan
      1 öronspottkörteln
      1 öronspottkörtlarna
      2 öronsus
      1 örontittare
      2 öronvärk
      2 öronvax
      1 orörda
      3 orörlig
      1 orörliga
      1 orörlighet
      1 orörligheten
      1 orörligt
      1 oroshärdar
      1 orostankar
      1 orpiment
    149 orsak
    265 orsaka
     90 orsakad
     67 orsakade
     14 orsakades
      8 orsakande
    280 orsakar
    299 orsakas
     30 orsakat
     19 orsakats
    221 orsaken
      1 orsakenorsakerna
    260 orsaker
     55 orsakerna
      1 orsakgrund
      2 orsaksfaktor
      1 orsaksfaktorer
      1 orsaksförhållande
      1 orsaksförhållandet
      1 orsaksmomenten
      3 orsakssamband
      1 orsakssambandet
      1 orsakssammanhang
      1 orsaksteori
      1 orsaksteorin
      1 orsakstyper
      2 örsnibben
      4 ort
     22 ört
      1 örtabok
      2 örtblad
      1 örtcigaretter
      7 orten
      2 örten
      2 Örten
      7 orter
     28 örter
      1 örterna
      1 örters
      1 orthokeratology
      1 orthokromatisk
      1 orthopedisk
      1 orthopoxvirus
      1 orthorexia
      2 orthos
      1 örtläkemedel
      1 örtmedicin
      3 örtmediciner
      1 örtmedicinska
      2 ortnamn
      3 orto
      4 ortodonti
      2 ortodontin
      5 ortodontisk
      1 ortodontiskt
      1 ortodontister
      3 ortodoxa
      1 ortodoxt
      1 ortofenylfenol
      2 ortogonalt
      8 ortografi
     10 ortografier
      1 ortografierna
      2 ortografin
      1 ortografiska
      1 ortohydroxiderivatet
      8 ortok
      2 ortomyxovirus
      1 ortopantomogram
      1 ortoped
      1 ortopeden
      1 ortopeder
      5 ortopedi
      3 ortopedin
      1 ortopedingenjörer
      7 ortopedisk
      1 ortopediska
      1 ortopediskt
      2 ortopné
      4 ortorektiker
      1 ortorektikers
      1 ortorektisk
      4 ortorektiska
     16 ortorexi
      1 ortorexia
      1 ortorombiska
      1 ortorombiskt
      8 ortos
      1 ortosbehandlingarna
      1 ortosen
      1 ortoser
      1 ortostatism
      1 örtstånd
      2 örtståndet
      1 örtterapier
      1 orubbade
      1 orvar
      2 orvietan
      1 orvieto
      5 os
      9 osa
      2 ösa
      6 osäker
      4 osäkerhet
      2 osäkerheten
      8 osäkert
      5 osäkra
      1 osaliga
      5 osammanhängande
      1 osanna
      3 osannolik
      2 osannolika
      5 osannolikt
      3 oscar
      1 oscarsgalan
      1 oscillationsfrekvens
      2 oscillerande
      1 oscillo
     22 oscilloskop
      1 oscilloskopbilden
      2 oscilloskopen
     13 oscilloskopet
      1 oscilloskopets
      2 osedligt
      1 osedvanligt
      1 oselektiva
      4 oseltamivir
      1 oserverats
      1 oshawa
      1 osiris
      1 osis
      1 osjälviska
      1 osjälvständig
      1 osjälvständigt
      1 oskadad
      2 oskadade
      1 oskadat
      1 oskadd
      2 oskadda
      1 oskadliga
      2 oskadliggöra
      1 oskadliggöras
      1 oskadliggörs
      1 oskar
      1 öskar
      1 osköljda
      1 oskrivna
      2 oskuld
      1 oskyddad
      5 oskyddade
      5 oskyddat
      1 oskyldig
      1 oskyldiga
      1 oskyldige
      1 osläckt
      5 osler
      1 oslo
      1 oslotrakten
      3 osmält
      2 osmältbara
      1 osmanska
      1 osme
      2 osmium
      1 osmo
      1 osmolaritet
      2 osmond
      2 osmoreglering
      5 osmos
      6 osmotisk
      2 osmotiska
      1 osmotiskt
      1 osorterad
      1 ospecificerade
      5 ospecifik
     15 ospecifika
      2 ospecifikt
      2 ospjälkade
     47 oss
      1 osseointegration
      1 osseointegrerade
      1 osseointegrering
      1 ossländerna
      1 osspelet
      6 ost
      1 öst
      4 Öst
      1 ostadiga
      2 ostadigheter
      1 ostadighetskänsla
      1 östafrikaner
      2 ostar
      2 östasiatiska
      3 Östasien
     10 osteit
      1 osteoartrit
      1 osteoklaster
      2 osteoklasterna
      1 osteoklasternas
      1 osteokondrodystropi
      1 osteokondros
      1 osteolys
      2 osteomalaci
      2 osteomyelit
      1 osteon
      1 osteopati
      3 osteopeni
      7 osteoporos
     20 osteosarkom
      1 osteoskelett
      1 osteotomi
      1 Österfärnebo
      2 Östergötland
      1 Östergötlands
      9 Österrike
      1 Österrikes
      1 Österrikeungern
      2 österrikisk
      3 österrikiska
      1 Österrikiska
      1 österrikiskamerikanske
      1 österrikiskbrittiska
      3 österrikiske
      1 österrikiskitalienska
      1 österrikiskungerske
      2 Östersjön
      1 Östersjöns
      1 Östersjösälarna
      4 Östersunds
      6 österut
      5 Östeuropa
      1 östeuropeiska
      1 Östgaard
      2 ostindien
      1 ostindisk
      3 östkusten
      2 östkustskolan
      3 östlig
      1 ostliknande
      1 östogenproduktionen
      1 ostört
      1 ostoyae
     19 östra
      3 Östra
     10 östradiol
      3 östriol
     68 östrogen
     10 Östrogen
      1 östrogena
      6 östrogenbehandling
      3 Östrogenbehandling
      2 östrogenberoende
     11 östrogener
      1 Östrogener
      1 östrogenerna
      2 Östrogenerna
     14 östrogenet
      8 Östrogenet
      5 östrogenets
      1 östrogenfasen
      1 östrogenfria
      1 östrogenfunktion
      1 östrogeninverkan
      1 östrogenkällor
      1 östrogenkörtlarna
      6 östrogennivåer
      9 östrogennivåerna
      1 Östrogennivåerna
      1 östrogenppiller
      1 Östrogenproduktion
      1 östrogenreceptor
      1 Östrogenreceptor
      6 östrogenreceptorer
      1 östrogenreceptorerna
      1 östrogenreceptormodulatorer
      1 östrogenreceptormodulerare
      2 östrogenreceptorn
      1 Östrogenreceptorn
      1 östrogenringar
      2 Östrogenringar
      1 östrogens
      1 östrogensyntes
      1 östrogent
      1 östrogentillförsel
      1 östrogenvärden
      1 östrogenverkan
      5 östron
      1 Östron
      1 östronet
      1 ostronskal
      1 ostsorter
      1 öststater
      1 Östsverige
      2 osunda
      1 osunt
     25 osv
      1 osymmetriska
      2 osynlig
      8 osynliga
      2 osynligt
      1 otäcka
      1 otakt
      3 otal
      1 otålbart
      4 otaliga
      1 otänkbart
      1 otäta
      1 otavit
      1 otestad
      1 other
      1 otherwise
      1 otidigt
      4 otillåtet
      3 otillåtna
      1 otillbörliga
      2 otillförlitliga
      1 otillfredsställande
      2 otillfredsställd
      1 otillfredsställda
      1 otillfredsställelse
      1 otillgängliga
     17 otillräcklig
      5 otillräckliga
     15 otillräckligt
      1 otit
      1 otites
      4 otitis
      1 otjänlig
      1 otoakustiska
      1 otolaryngolog
      1 otorhinolaryngologi
      3 otoskop
      4 otoskopet
      2 otpf
      2 otränad
      1 otränade
      1 otrevlig
      1 otrevligheter
      1 otrevligt
      1 otrogen
      1 otrohet
      1 otroheten
      1 otrolig
      3 otroligt
      2 otrygg
      1 otrygga
      2 otryggambivalent
      1 otryggdesorganiserad
      2 otryggundvikande
      2 otsj
      1 otsuka
      6 otto
      1 otukt
      1 otur
      1 oturen
      2 otvetydiga
      1 otvivelaktligen
      2 otydlig
      4 otydliga
      1 otydligare
      1 otympliga
      4 otypiska
      2 otypiskt
     13 Ötzi
      5 Ötzis
      1 Ötztalalperna
      1 oumbärlig
      2 ounce
      2 oundviklig
      1 oundvikliga
      1 oundvikligt
      1 oupphettade
      2 oupphörligen
      1 oupplösligen
      1 oupplysta
      2 ouppmärksam
      4 ouppmärksamhet
      1 ouppmärksammade
      2 oupptäckta
      1 our
      1 ourselves
      2 out
      1 outbildad
      1 outhärdlig
      1 outhärdliga
      1 outhärdligt
      2 output
      1 outsläcklig
      1 outspjälkad
      1 ouwens
      5 öva
      4 ovaccinerade
      1 oväder
      2 oval
      9 ovala
      3 ovale
      1 ovalformade
      1 ovalutionssmärta
     37 ovan
      3 ovana
      1 ovandelen
     30 ovanför
      1 ovanifrån
      1 ovanirån
      2 ovanjordiska
      1 ovanjordiskt
      1 ovanjordsdelen
     59 ovanlig
     48 ovanliga
     19 ovanligare
      3 ovanligaste
      1 ovanliggande
    117 ovanligt
      1 ovanligtbr
      1 ovannämnda
      1 ovanor
     13 ovanpå
      6 ovansida
      8 ovansidan
      2 ovansjö
     13 ovanstående
      3 oväntad
      2 oväntade
      1 oväntat
      1 övar
      1 ovarial
      2 ovarialcancer
      3 ovarialsvikt
      2 ovarialtorsion
      3 ovariell
      1 ovarier
      1 ovarierna
      7 ovariesyndrom
      1 ovariet
      1 ovarii
      3 ovariotomi
      2 ovariotomier
      4 ovariotomin
      1 ovariotomins
      1 ovariotomist
      2 ovarium
      2 övärlden
      2 övas
      2 oväsen
      1 oväsentlig
      1 ove
      1 övegripande
      1 oven
    666 över
     12 Över
      7 överaktiv
      2 överaktiva
      1 överaktiverad
      1 Överaktiveringen
      2 överaktivitet
      1 överaktivitetssymtom
      1 överaktivt
     16 överallt
      2 överansträngd
      1 Överansträngd
      1 överansträngda
     11 överansträngning
      1 överansträngningen
      1 överanvänder
      1 överanvändning
      1 överanvänts
      1 överarmen
      2 överarmens
      3 överarmsbenet
      1 överbebodd
      1 överbefolkad
      1 överbefolkning
      2 överbelastar
      1 överbelastas
     10 överbelastning
      1 Överbelastning
      2 överbeskyddande
      2 överbevisad
      1 överbevisats
      3 överblick
      1 överblicka
      1 överblickas
      1 överbliven
      2 överblivna
      2 överdel
      1 överdelar
      1 överdelsfri
      1 överdiagnostiserad
      1 Överdiagnostisering
      1 överdirektion
      1 överdirektör
      8 överdos
      2 Överdos
      2 överdoser
      2 överdosera
      1 överdoserar
      5 överdosering
      1 överdra
      1 överdragen
      1 överdrift
      2 överdriva
     20 överdriven
      1 Överdriven
     12 överdrivet
      7 överdrivna
      1 Överdrivna
     18 överens
      1 överenskommas
      1 överenskommelser
      2 överensstämma
      1 överensstämmande
      3 överensstämmelse
      1 överensstämmelsen
     14 överensstämmer
      1 överfallen
      1 överfamilj
      5 överflöd
      2 överflödig
      3 överflödiga
      1 överflödigt
      1 överflyglades
      2 överflyttades
      1 överflyttas
     11 överför
     14 överföra
      1 överförandet
     28 överföras
      7 överförbar
     13 överförbara
      1 överförbart
      3 överförd
      4 överförda
      1 överförde
     10 överfördes
      1 överförfriskade
     21 överföring
      8 Överföring
      4 överföringar
      2 överföringarna
      7 överföringen
      1 Överföringen
      1 överföringsfrekvensen
      1 överföringsrör
      2 överföringsrören
      2 överföringssätt
      1 överföringsvägen
     46 överförs
      2 överfört
      6 överförts
      1 överfulla
     19 övergå
     23 övergående
      1 Övergående
      6 övergång
      1 Övergång
      1 övergångar
      7 övergången
      3 Övergången
      2 övergångsåldern
      1 övergångsbesvär
      2 övergångsepitelcancer
      1 Övergångsepitelcancer
      1 övergångsperiod
      1 övergångsperioden
      5 övergångsställe
      1 Övergångsställe
      5 övergångsställen
      1 övergångsställets
      1 övergångstid
      1 övergångstillstånd
     26 övergår
      7 övergått
      1 övergavs
      3 överge
      1 överges
      1 övergetts
      5 övergick
      1 övergivande
      1 övergivit
      2 övergivits
      3 övergivna
      1 övergödning
      6 övergrepp
      1 Övergrepp
     11 övergripande
      2 Övergripande
      1 Övergripligt
      3 överhanden
      2 överhängande
      1 överhettas
      1 överhettning
      1 överhöljda
      1 överhud
      1 Överhud
      5 överhuden
      1 Överhuden
     11 överhuvudtaget
      1 överinformation
      1 överinlärda
      1 överinlärning
      1 överinseende
      1 överintelligens
      4 överjaget
      1 överkäke
      3 överkäken
      7 överkänslig
      6 överkänsliga
     34 överkänslighet
      6 Överkänslighet
      1 Överkänsligheten
      5 överkänslighetsreaktion
      8 överkänslighetsreaktioner
      2 överkänslighetssymtom
      1 överkapacitet
      1 överklaga
      1 överklagades
      1 överklagan
      1 överklagas
      6 överklassen
      2 overklig
      3 overkliga
      1 overklighet
      2 overklighetskänsla
      4 overklighetskänslor
      1 overklighetskänslorna
      2 overkligt
      1 överkomlig
      2 överkomma
      4 överkonsumtion
      2 Överkonsumtion
      5 överkropp
      2 överkroppen
      1 overksam
      1 overksamma
      1 overksamt
      1 överkuporna
      2 överlack
      1 överlag
      1 överläggs
      1 överlagrad
      2 överlagras
      1 överlagrats
      1 överlagringseffekter
      3 överlägsen
      2 överlägsenhet
      4 överlägset
      1 överlägsna
      3 överläkare
      2 överläkaren
      2 överlämna
      1 överlämnades
      1 överlämnande
      1 överlämnar
      1 överlapp
      1 överlappande
      1 overlappar
      5 överlappar
      2 överläppen
      1 Överläppen
      1 överlappning
      1 Överlappningen
      2 överlåtas
      1 överledningen
     31 överleva
      7 överlevande
      1 Överlevanden
      9 överlevde
     26 överlever
     29 överlevnad
      5 överlevnaden
      1 Överlevnaden
      1 överlevnadicke
      1 överlevnadsångest
      3 överlevnadschansen
      1 överlevnadschanserna
      1 överlevnadsdriften
      2 Överlevnadsfrekvensen
      1 överlevnadsinstinkt
      1 överlevnadsmål
      2 överlevnadsmöjligheter
      1 överlevnadsstatistiken
      1 överlevnadsstrategi
      2 överlevnadstid
      2 överlevnadstiden
      1 Överlevnadstiden
     13 överlevt
      1 överlista
      2 övermäktiga
      1 övermäktigt
      1 övermanna
      1 övermänsklig
      1 övermänskliga
      1 övermaskuliniserad
      1 övermättnaden
      3 övernaturlig
      8 övernaturliga
      1 övernaturligas
      5 övernaturligt
      1 övernormalt
      1 Överoptimism
      1 överoptimistiska
      1 överordnade
      2 överordnat
      2 överproduceras
      2 överproduktion
      1 Överproduktion
      1 överpronation
      3 överraskade
      4 överraskande
      1 överraskat
      1 överraskats
      2 överraskning
      1 överraskningar
      2 överreagerande
      1 överreagerar
      3 överreaktion
      1 överreaktioner
      2 överrepresentation
      4 överrepresenterade
      1 överrepresenterat
      1 överrinningsinkontinens
      1 överrock
      1 överrörlighet
      1 överrörlighetssyndrom
      1 överröstas
      1 övers
      9 översatt
      1 Översatt
      5 översättas
      1 översatte
      2 översätter
      1 översattes
      6 översättning
      1 översättningar
      2 översättningen
      1 översatts
      3 översätts
      1 översekretion
      1 översignalering
     10 översikt
      2 Översikt
      1 Översikten
      1 översikter
      1 översiktlig
      1 Översiktlig
      1 Översjälen
      1 Överskådligt
      2 överskatta
      2 överskattar
      1 överskattas
      8 överskott
      4 överskottet
      1 Överskottet
      1 överskottsfett
      4 överskottshud
      1 överskottslager
      1 överskottsslam
      1 överskottsslamet
      1 överskottsvärmen
      2 överskottsvätska
      5 överskrida
      1 överskridas
      6 överskrider
      1 överskridit
      1 överskrids
      1 överskuggande
      7 överst
      1 Överst
      6 översta
      2 överstatliga
      1 översteg
      1 överstelöjtnant
      2 överstiga
     17 överstiger
      1 överstigt
      1 överstimulera
      1 överstimuleras
      1 överstimulering
      2 översträckning
      1 översträcks
      1 överstyr
      1 Överstyrelsen
      4 översvämningar
      1 översvämningsområde
      2 översyn
      1 översynthet
      1 Översynthet
      3 överta
      1 övertag
      1 övertagande
      1 övertaget
      1 övertagit
      2 övertaliga
      1 övertandläkare
      1 övertog
      2 övertogs
      2 övertoner
      1 övertonsrik
      1 överträda
      1 överträdas
      1 överträdelser
      1 överträffande
      1 överträffar
      1 överträning
      9 övertryck
      1 Övertryck
      3 övertrycksandning
      1 övertrycksmiljö
      1 övertrycksventilation
      2 övertyga
      5 övertygad
      4 övertygade
      4 övertygande
      1 övertygas
      2 övertygelse
      1 överväg
      7 överväga
     10 övervägande
      7 övervägas
      5 överväger
      1 övervägs
      5 övervaka
      3 övervakad
      1 övervakade
      1 övervakades
      2 övervakande
      9 övervakar
     10 övervakas
      1 övervakat
     25 övervakning
      2 Övervakning
      4 övervakningen
      1 Övervakningen
      1 övervakningsdatorer
      1 övervakningsmål
      3 överväldigande
      1 övervåningen
      2 övervätskning
      3 överväxt
     33 övervikt
      2 Övervikt
      1 övervikten
      2 överviktig
     15 överviktiga
      1 Överviktigas
      1 överviktigt
      1 övervinna
      1 övervinner
      1 övervintra
      1 övervintrande
      4 övervintrar
      1 övervintringsknopparna
      1 ovetandes
      1 ovidius
      1 oviktigt
      1 ovilja
      1 oviljan
      1 ovillig
      3 ovilliga
      1 ovipar
      1 oviss
      1 övning
     12 övningar
      1 övningarna
      1 övningen
      2 ovocyst
      1 ovocyten
     94 övre
      4 Övre
      5 övrig
      4 Övrig
    111 övriga
     15 Övriga
     39 övrigt
      8 Övrigt
      1 ovulation
      1 ovulationen
      1 ovulerade
      2 owen
      1 own
      1 ox
      1 oxacillin
      1 oxalacetat
      1 oxalat
      1 oxalater
      1 oxalsyra
      3 oxar
      1 oxazepam
      1 oxbär
      1 oxcytocin
      3 oxford
      1 oxforduniversitetet
      2 oxgalla
      1 oxhuvuden
      3 oxid
      1 oxidas
     15 oxidation
      1 oxidationen
      3 oxidationsmedel
      1 oxidationsmedlet
      1 oxidationsprodukt
      1 oxidationstal
      2 oxidativ
      1 oxidativa
      1 oxidativt
      1 oxidator
      1 oxider
      3 oxidera
      1 oxiderade
      1 oxiderades
      8 oxiderande
      6 oxiderar
     11 oxideras
      4 oxiderat
      1 oxidering
      1 oxideringsämnen
      1 oxidopamin
      1 oxihemoglobin
      1 oxiketoner
      1 oxitetracyklin
      4 oxygen
      1 oxygenol
      1 oxyhemoglobin
     47 oxytocin
      1 oxytocinaktivitet
      1 oxytocinaktiviteten
      6 oxytocinet
      2 oxytocinnivåerna
      3 oxytocinreceptorer
      1 oxytocinutsöndring
      5 oxyuranus
      1 ozein
     15 ozon
      1 ozonbehandling
      2 ozonet
      1 ozonhål
      2 ozonhålet
      1 ozonhalten
      3 ozonlagret
      1 ozonmolekylerna
      1 ozonnerbrytande
      1 ozonpåverkande
      1 ozontekniken
     34 p
      1 [p]
      2 pa
   8067 på
      1 [pa�a]
      1 påbjuds
      1 pablo
      6 påbörja
      5 påbörjad
      3 påbörjade
      4 påbörjades
      1 påbörjandet
      5 påbörjar
     21 påbörjas
      3 påbörjat
      4 påbörjats
      1 påbyggnadsår
      1 påbyggnadskurser
      4 påbyggnadsutbildning
      1 påbyggnadsutbildningar
      8 pacemaker
      1 pacificera
      1 pacifistisk
      1 pacifistiskt
      3 packa
      1 packad
      2 packade
      2 packas
      2 packningar
      1 packningen
      1 packsten
      2 paco
      6 pacs
      1 pacset
      2 padar
      1 padda
      2 pådrivande
      1 påengelska
      1 påfallade
      7 påfallande
     10 påföljande
      1 påföljd
      1 påföljden
      1 påföljder
      2 påfresta
      7 påfrestande
      4 påfrestning
     16 påfrestningar
      1 påfrestningen
      1 påfunnits
      1 påfyllnad
      5 påfyllnadsdos
      2 påfyllning
     10 pågå
     16 pågående
      1 pågar
     39 pågår
      8 pågått
      1 page
      2 paget
      1 pagets
      7 pågick
      1 påhittad
      1 påhittade
      1 påhittat
      1 paideia
      1 paiderastia
      1 paidos
      2 pain
      2 pais
      1 påkalla
      1 påkallar
      1 påkallats
      3 paket
      1 paketering
      1 paketet
      1 pakethållaren
      6 pakistan
      4 paklitaxel
      1 påkommande
      2 påkommen
      1 påkomna
      1 påkörd
      1 påkörningar
      1 pakter
      1 pal
      2 pålägg
      1 påläggning
      1 palaquium
      1 pålästa
      1 palatoglossus
      1 palats
      1 palb
      1 palditaxol
      1 paleoantropologerna
      3 paleolitikum
      2 paleolitisk
      3 paleolitiska
      1 paleontologen
      1 palestinska
      1 paletter
      5 palilali
      1 palilalia
      1 palilalie
      1 pålimmade
      2 pálin
      2 pålitlig
      5 pålitliga
      2 pålitligare
      1 pålitligaste
      1 pålitlighet
      2 pålitligt
      1 pallescens
      6 palliativ
     21 pallidum
      1 pallidumspecifika
      1 palmarerytem
      1 palme
      4 palmer
      1 palmerister
      2 palmers
      1 palmitinsyra
      1 palmolivepeet
      1 palmolivetvålen
      4 palmolja
      5 palpation
      1 palpera
      1 palperbar
      1 palpering
      5 palpitationer
      3 pålrot
      6 päls
      1 pälsar
      1 pälsbyxor
      1 pälsbyxorna
      3 pälsdjur
      1 pälsdjuret
      1 pälsdjursallergi
      6 pälsen
      1 pälshandlare
      1 pälslösa
      1 pälsprodukter
      1 pälsrock
      1 pälssorter
      2 paltkoma
      1 paltschwimen
      1 palynologi
      1 påmålning
      1 pamela
      1 pamflett
      2 påmind
      3 påminde
      3 påminna
      1 påminnande
     35 påminner
      1 påmint
      1 pamp
      1 pampig
      3 panama
      3 panamic
      1 panchakarma
      1 pancicii
      1 pancoasttumörer
      5 pancreas
      1 pancreasgången
      4 pancreaticus
      1 pancres
      8 pandas
      1 pandaskriterierna
      1 pandasundergrupp
     11 pandemi
      1 pandemia
      8 pandemier
      2 pandemierna
      2 pandemin
      2 pandemisk
      1 pandemiskt
     10 pandemrix
      1 pandemrixutlöst
      1 paneler
      1 panencefalit
     11 panik
     18 panikångest
      1 panikångesten
      1 panikartad
      5 panikattack
     12 panikattacker
      1 panikkänslor
      1 paniksituation
      8 paniksyndrom
      5 pankreas
      2 pankreassaft
      1 pankreassaften
      7 pankreatit
      2 pankuroniumbromid
      3 panna
      4 pannan
      1 pannbenet
      1 pannbenets
      1 pannloben
      1 pannlobens
      1 pannlobsdemens
      1 pannonicus
      1 pannor
      1 pannrum
      5 pannsten
      1 pannstensbildande
      2 panocod
      3 pans
      4 panss
      1 panterfläckig
      5 panterflugsvamp
      1 pantermusseron
      1 pantermusseronen
      1 pantherina
      1 pantoprazol
      1 pantotensyra
      1 pånyttfödas
      1 panzona
      1 pao
      3 paolo
      1 papatasii
      1 papaverin
      1 papegojfåglar
      1 papegojor
      2 papegojsjuka
      1 papegojsjukan
      2 påpeka
      2 påpekade
      1 påpekades
      6 påpekar
      1 påpekas
      2 påpekat
      1 papel
      1 papers
      3 papilla
      7 papillae
      3 papillär
      1 papillarmuskler
      2 papillärt
      1 papiller
      1 papillnekros
      5 papillomavirus
      1 papillomvirus
      1 papillösa
      2 papler
      1 papp
      2 pappa
      1 pappaersaktig
      1 pappan
     15 papper
      5 papperet
      1 papperets
      2 pappers
      1 pappersdokument
      1 pappersfibrer
      1 pappersförpackningar
      3 pappershanddukar
      2 pappershandduken
      1 pappersida
      1 pappersindustri
      1 papperskorgar
      1 papperskromatografi
      2 papperslapp
      1 papperslappar
      1 pappersmaskinerna
      4 pappersmassa
      1 pappersmassor
      1 papperspåse
      1 papperspositiv
      2 pappersremsa
      1 pappersremsan
      1 pappersservetter
      1 papperstunna
      1 pappersutskrift
      1 papphylsa
      1 pappmaskin
      1 pappografi
      1 pappren
      3 pappret
      1 papprullen
      1 papsmear
      3 papua
      1 papules
      2 papyri
      7 papyrus
      1 papyrusen
      1 papyrusfoster
      2 papyrusrullar
      1 papyrusrullen
    105 par
      1 pär
      7 para
      3 paraaminosalicylsyra
      1 paracaskulturen
      1 paracellulär
      1 paracellulära
      1 paracelsism
     11 paracelsus
     10 paracetamol
      1 parad
      1 parade
      1 paradigm
      1 paradigmet
      2 paradigmskifte
      1 paradisartade
      1 paradise
      5 paradiset
      1 paradox
      3 paradoxal
      1 paradoxala
      3 paradoxalt
      1 paradoxus
      1 paraduniform
      1 parafasi
      1 parafasier
      1 parafernalia
      1 parafila
      9 parafili
      9 parafilier
      2 parafilierna
      3 parafilin
      2 parafimos
      1 parafollikullära
      1 paraföreningar
      2 parafyletisk
      1 paragonimiasis
      1 paragonimus
      1 paraguayensis
      1 parainfluensa
      2 parainfluensavirus
      1 parainfluensvirus
      2 parakeratos
      1 parakresol
      1 parakrin
      1 parakusi
      1 parallell
      9 parallella
      1 paralleller
     13 parallellt
      1 paralympics
      2 paralys
      3 paralysera
      2 paralyserar
      2 paralytica
      1 paralytisk
      2 paramatma
      1 paramedicin
      1 paramedicinen
      1 paramenstruell
      3 parametern
     10 parametrar
      2 parametrarna
      1 paramilitära
      1 paraminobensoesyra
      2 paraminobensoesyran
      1 paraminobensoesyrans
      1 paramyxoviridae
      1 paramyxovirus
      1 paranensis
      1 paraneoplastiska
      1 paraneoplastiskt
     19 paranoia
      1 paranoian
      1 paranoianätverket
     19 paranoid
      6 paranoida
      1 paranoide
      1 paranötter
      3 paraorange
      3 parapares
      3 parapertussis
      1 parapertussisstammar
      1 paraphimosis
      2 paraplegi
      1 paraplegiker
      1 paraplybeteckning
      2 paraplyterm
      1 parapneumonisk
      1 paraprotein
      1 paraproteinemi
      2 paraproteiner
      1 paraproteinet
      1 parapsykologin
      1 parapsykologisk
      4 parar
      1 paras
     10 parasit
      1 parasitangrepp
      1 parasitära
      1 parasitcystor
     35 parasiten
      2 parasitens
     36 parasiter
      2 parasitera
      9 parasiterande
      8 parasiterar
     13 parasiterna
      1 parasitinfektion
      1 parasitinfektioner
      5 parasitisk
      5 parasitiska
      1 parasitismen
      2 parasitmask
      3 parasitmasken
      1 parasitologi
      1 parasitología
      4 parasitsjukdom
      1 parasitsjukdomar
      1 parasitsjukdomen
      1 parasitspecifika
      1 parasitsvampar
      3 parasomni
      3 parasomnier
      2 parasomnierna
      4 parasympatiska
      1 parat
      1 paratetrapares
      1 paratyroidea
      1 paratyroideahormon
      2 paratyroideahormonet
      1 paraventrikulära
      5 parbildning
      3 parbladiga
      2 parc
      1 parcopresis
      1 pardelade
      1 pardinum
      2 paré
      1 parenkymliknande
      1 parent
      1 parentchild
      2 parenteral
      1 parenterala
      1 parenteralt
      3 parentes
      7 pares
      1 pareser
      4 parestesi
      2 parestesier
      4 paret
      1 parflikiga
      7 parfym
      5 parfymämnen
      1 parfymburkar
      2 parfymer
      1 parfymera
      1 parfymerades
      1 parfymerat
      1 parfymering
      1 parfymfri
      1 parfymfria
      1 parfymkulor
      1 parfymtillverkning
      1 pariboy
      1 parietal
      1 parietala
      3 parietalceller
      2 parietalcellerna
      8 parietalloben
      2 parietallobslesioner
      1 parietoccipitallobotomi
      1 parig
      3 pariga
     30 paris
      1 parisbesök
      1 parisergrönt
      1 parisgrönt
      1 parisiska
      2 parissyndromet
      1 paritalloben
      3 park
      4 parker
      1 parkera
      1 parkeringshus
      1 parkeringsläge
      1 parkeringsövervakning
      2 parkinson
      2 parkinsonism
      1 parkinsonliknande
      1 parkinsonpatienter
     18 parkinsons
      1 parkki
      1 parklandsformel
      1 parkmiljöer
      1 parkträd
      1 pärla
      1 parlament
      1 parlamentariska
      2 parlamentet
      1 pärldykare
      1 pärlliknande
      3 pärlor
      1 pärlring
      1 parlys
      8 parning
     13 parningen
      1 parningens
      1 parningsberedskapen
      1 parningsbeteende
      1 parningsdräkt
      1 parningsinriktade
      2 parningslekar
      3 parningsorgan
      1 parningsorganen
      1 parningssäsongen
      1 parningstiden
      1 parodii
      1 parodontal
      1 parodontala
     12 parodontit
      1 parodontiten
      1 parodontolog
      2 parodontologi
      1 päron
      2 päronformad
      2 päronpest
      1 päronträd
      1 parosmi
      1 parotiskörteln
      1 parotiskörtelns
      2 parotit
      1 parotitvirus
      4 parotitviruset
      1 parövningar
      1 paroxetin
      1 paroxysm
      1 paroxysmal
      1 paroxysmós
      1 parr
      1 parrs
      3 pars
      3 parsamtal
      5 part
      4 parten
     10 partenogenes
      1 partenogeneshandling
      2 partenogenetiskt
      1 partens
      3 parter
      3 parti
      1 partialdrift
     12 partialtryck
      7 partialtrycket
      1 particle
     18 partiell
      6 partiella
      4 partiellt
      2 partier
      1 partierna
      1 partihandel
      2 partikel
      1 partikelaccelerator
      1 partikelacceleratorer
      1 partikelenergi
      1 partikelfysik
      1 partikelhalt
      1 partikeln
      1 partikelslag
      2 partikelstrålning
     21 partiklar
     10 partiklarna
      3 partiklarnas
      1 partiklars
      1 partiska
     33 partner
      1 partnerbrev
      9 partnern
      1 partnerns
      1 partnerrelationer
      6 partners
      1 partnership
      3 partnerskap
      1 partre
      1 pärts
      1 partum
      2 partus
      1 partydrog
      6 paruresis
      1 parvifolius
      1 parvis
      6 parvovirus
      1 parvum
     28 pas
      1 [pas]
      6 påsar
      2 påsarna
      1 pasbehandling
      1 pasbehandlingen
      1 påsbyten
      3 påsdialys
      4 påse
      3 påsen
      1 pasi
      1 påsk
      1 påsketeje
      1 påsketet
      2 påsklilja
      2 påskliljan
      1 påskliljans
      1 påskliljor
      1 påskön
      5 påskynda
      1 påskyndad
      6 påskyndar
      1 påskyndas
      2 påslag
      2 påslaget
      1 påslagna
     24 pass
     12 passa
      2 passade
     14 passage
      1 passagemetabolism
      3 passagen
      1 passagerarflygplan
      1 passagerarna
      1 passageväg
      4 passande
     23 passar
     35 passera
      1 passerande
     39 passerar
     13 passerat
      1 passerats
      2 passet
      2 passform
      1 passformen
      1 passion
      1 passitometoden
     11 passiv
      3 passiva
      1 passivaggressiv
      1 passivisera
      3 passivitet
     10 passivt
     27 påssjuka
      1 påssjukans
      1 påssjukedelen
      1 påssjukemeningit
      2 påssjukevirus
      3 passtreptomycin
      3 pasta
      2 påstå
      2 påstådd
      7 påstådda
      3 påstående
     16 påståenden
      1 påståendena
      3 påståendet
      1 pastaform
      1 pastan
      9 påstår
     18 påstås
      3 påstått
      5 påståtts
      1 pastell
      1 pastellfärg
      2 pasteur
      1 pasteurella
      1 pasteurinstitutet
      1 pastiller
      5 påstod
      3 påstods
      1 pastor
      1 pastöriseringen
      1 pastöriseringsprocessen
      1 påtäffades
     11 påtaglig
      6 påtagliga
      1 påtagligare
      1 påtagligast
     11 påtagligt
      2 påtalar
      1 påtalats
      2 patanjali
      1 patanjalis
      4 pataus
      1 patéer
      1 pateientens
      1 patellaluxation
      1 patellarreflex
     11 patent
      2 patenterad
      1 patenterade
      2 patenterades
      2 patentet
      1 patentmedicin
      1 patentmediciner
      1 patentmedicinerna
      1 patentskyddade
      1 patenttid
      1 paterson
      1 pathogenesis
      1 pathologica
      3 pathological
      2 pathos
      1 páthos
      1 pathway
      1 pati
     72 patient
      2 patientdata
      2 patientdatalagen
      1 patientdrivna
    387 patienten
      1 patientenförsökspersonen
      1 patientenklienten
     96 patientens
      1 patientensföräldrarnas
      2 patientensförsökspersonens
      2 patientensklientens
      1 patientent
    323 patienter
      1 patienterkälla
     74 patienterna
      3 patienternas
      2 patientfall
      1 patientfallens
      1 patientfokus
      1 patientföljsamhet
      1 patientföreningen
      4 patientgrupp
      5 patientgruppen
      7 patientgrupper
      1 patientgrupperna
      1 patientinformationleaflet
      1 patientinformationsblad
      6 patientjournal
      1 patientjournaler
      1 patientjournallagen
      1 patientklientel
      1 patientläkarerelationen
      1 patientlift
      3 patientlyft
      3 patientlyftar
      1 patientlyftens
      1 patientnära
      1 patientöversikten
      1 patientprover
      1 patientrelaterade
      7 patients
      1 patientsäkerhet
      4 patientsäkerhetslagen
      1 patientstöd
      1 patientsystem
      1 patientunderlag
      1 patientutbildning
      1 patientvård
      1 patiet
      1 patietens
     10 patofysiologi
      1 patofysiologin
      2 patofysiologisk
     14 patogen
     12 patogena
      1 patogenen
      4 patogener
      2 patogenerna
      8 patogenes
      1 patogenet
      2 patogenets
      1 patogengruppen
      1 patogenicitet
      2 patogenitet
      3 patogent
      1 patognomona
      2 patognomont
     14 patologi
      2 patologin
      1 patologins
      1 patologisera
      8 patologisk
     22 patologiska
      1 patologiskanatomisk
      8 patologiskt
      1 patos
      7 påträffades
     22 påträffas
     11 påträffats
      1 påträngande
      1 patria
      1 patriarken
      1 patricio
      4 patrick
      1 patroner
      1 patronformat
      1 patrull
      1 patrullerande
      1 patrulleringsverksamhet
      1 påtryckning
      2 påtryckningar
      1 patt
      1 patta
      1 pattabhi
      1 pattern
      1 patterns
      2 påtvinga
      2 påtvingad
      1 påtvingas
      1 påtvingat
      3 paucibacillär
      1 pauciflorus
      1 pauksch
     15 paul
      1 paulescu
      3 pauser
      1 pausering
      1 pauseringsmönster
      1 pauseringstid
      1 påväxt
      1 påve
      1 påvebulla
      3 pavel
      3 påven
      1 påvens
    105 påverka
      7 påverkad
     29 påverkade
      3 påverkades
    105 påverkan
      2 påverkande
      1 påverkansgrad
      1 påverkansområden
    226 påverkar
    116 påverkas
      7 påverkat
      2 påverkats
      1 påverkningar
      1 påverks
      1 påvestaden
     36 påvisa
      2 påvisad
      7 påvisade
      5 påvisades
     13 påvisar
     23 påvisas
      5 påvisat
     18 påvisats
      3 påvisbar
      5 påvisbara
      1 påvisbart
      3 påvisning
      2 pavlov
      1 pavor
      1 pavulon
      1 paxillus
      1 paxton
      1 pb
      1 pbo
      4 pbp
      1 pbproteinerna
      2 pc
      1 pcantikropparna
      4 pcb
      1 pci
      1 pcinstickskort
      1 pcit
      1 pclr
      3 pco
      1 pcos
      3 pcp
     15 pcr
      1 pcrdetektion
      1 pcrdiagnostiken
      1 pcrprodukt
      2 pct
      1 pcv
      1 pd
      2 pdator
      7 pdatorer
      1 pdatorerna
      5 pdatorn
      1 pdv
      2 pe
      3 peak
      1 peakday
      1 peakflowmeter
      1 péan
      1 peang
      2 peanger
      1 péans
      1 pearce
      6 pearl
      6 pearlindex
      1 pechbländets
      1 pectinata
      3 pectoris
      3 pectus
      1 peczlsy
      1 peczly
      1 pedagog
      1 pedagogen
      2 pedagogik
      1 pedagogiken
      5 pedagogisk
      6 pedagogiska
      4 pedagogiskt
      1 pedaldriven
      1 pedalrörelser
      1 pedanius
      1 pederast
      1 pederaster
      1 pederastförhållanden
     12 pederasti
      7 pederastiförhållanden
      8 pederastin
      1 pederastisk
      2 pederastiska
      1 pederastiskt
      2 pedersen
      1 pediater
      2 pediatric
      2 pediatrics
      5 pediatrik
      1 pediatriker
      4 pediatrisk
      4 pedikyr
      5 pedis
      1 pedodonti
      1 pedofil
      1 pedofili
      1 pedriatriken
      1 peelande
      2 peeling
      2 peelingeffekt
      4 peep
      2 peer
      1 peet
      3 pef
      3 peg
      1 pegen
      2 pehr
      1 pek
      2 peka
      1 pekannötter
     28 pekar
      5 pekat
      1 pekfingrar
      1 pekskärmstelefon
      1 pel
      2 pelele
      1 peligot
      1 pelle
      1 pellets
     14 pellucida
      1 pelviotomi
      1 pelvospondylit
      1 pemfigoid
      2 pemolin
      1 pemphigus
      1 pencillin
      1 pencillinerna
      1 pendelrörelser
      1 pendeltåg
      1 pendla
      2 pendlar
      1 pendlat
      3 penetration
      1 penetrationssex
      5 penetrera
      1 penetrerade
      3 penetrerar
      3 penetreras
      2 penetrerat
      1 penetrerats
      1 penetrering
      1 penfieldkanadensare
     20 pengar
     45 penicillin
      2 penicillinallergi
      1 penicillinallergier
      1 penicillinas
      1 penicillinaset
      2 penicillinbehandling
      1 penicillinbindande
      5 penicilliner
      2 penicillinet
      4 penicillininbindande
      1 penicillinkänsliga
      1 penicillinproduktionen
      1 penicillinresistens
      2 penicillium
     72 penis
      1 penisavund
      1 penisbasblockad
      2 penisben
      2 peniscancer
      7 penisen
      1 penisens
      2 penisförstoring
      2 penisfraktur
      1 penisprotes
      2 penisroten
      2 penisskaftet
      1 penistillväxten
      1 penisvävnaden
      1 penna
      1 pennor
      2 pennsylvania
      1 pensée
      1 pensel
      1 penselformigt
      2 penselmögel
      1 pension
      1 pensionärer
      2 pensionerades
      1 penslas
      1 pentaploid
      1 pentasa
      1 pentothal
      1 pentrerande
      2 people
      1 peplus
      1 pepo
      1 pepparmint
      1 pepparmynta
      1 pepprigt
      1 pepsi
      3 pepsin
      4 pepsinogen
      1 peptid
      1 peptidas
      1 peptidbryggor
      1 peptiden
      9 peptider
      5 peptiderna
      6 peptidhormon
      3 peptidhormoner
      5 peptidkedja
      2 peptidkedjan
      2 peptidkedjor
      1 peptidlänkar
      1 peptidlösning
      1 pepys
    269 per
      1 peramivir
      6 perättiksyra
      2 perce
      2 percentilen
      1 percentiler
     12 perception
      6 perceptionen
      1 perceptioner
      1 perceptions
      1 perceptionsfunktionerna
      1 perceptionsstörning
      2 perceptuell
      1 percutan
      1 peredo
      2 perenna
      1 perennis
      2 peres
      1 peretto
      1 perez
      1 perfect
      8 perfekt
      3 perfekta
      1 perfektionism
      1 perforerad
      1 perforerade
      1 perforeras
      1 perforering
      1 perforeringar
      5 performance
      3 perfringens
      1 perfuserar
      1 perfusion
      1 perfusionist
      3 perfusionisten
      1 perfusionistens
      3 perfusionister
      1 perfusionistkåren
      1 perfusionistutbildning
      1 perfusionstrycket
      1 pergolid
      2 perianal
      1 periarterit
      1 periartrit
      6 pericyter
      1 perietal
      9 perifer
     44 perifera
      1 periferala
      1 periferiseendet
      8 perifert
      1 perifornikala
      1 perihilära
      1 perikard
      2 perikardiet
      6 perikardit
      1 perikardium
      1 perinatal
      1 perinatala
      1 perineum
     64 period
      1 periodare
     20 perioden
     39 perioder
      4 perioderna
      1 periodicitet
      1 periodiciteten
      1 periodicitetsanalys
      1 periodicitetsteorin
      4 periodisk
      2 periodiska
      2 periodiskt
      1 periodontologi
      1 periodprevalens
      3 periodvis
      2 periostit
      1 peripneumoni
      1 peristaltik
      6 peristaltiken
      7 peristaltiska
      1 perithecium
     11 peritonealdialys
      3 peritoneum
      4 peritonit
      1 perkin
      1 perkloretylen
      1 perkussion
      3 perkutan
      1 perlane
      1 perlino
      1 perlman
      4 perls
     44 permanent
      9 permanenta
      1 permeabel
      1 permeabelt
      4 permeabilitet
      1 permeabiliteten
      1 permetrin
      1 permissionsuniform
      2 perniciös
      1 peroneuspares
      7 peroralt
      1 peroxid
      1 peroxidas
      1 peroxidaser
      1 peroxider
      1 peroxidfamiljen
      1 perpetuell
      1 perrektalt
      1 perrier
      1 perserna
      1 perseveratio
      2 perseveration
      1 perseverationer
      1 perseverativa
      1 persevero
      2 persicum
      2 persien
      1 persikaplommonkörsbärmandel
      2 persilja
      1 persisk
      4 persiska
      1 persiskt
      1 persistent
      1 persistenta
      2 persisterande
      1 persoenr
    393 person
      1 persona
     43 personal
      2 personaladministration
      1 personalbrist
     13 personalen
      2 personalens
      1 personalfrånvaro
      1 personalinvesteringar
      1 personalkostnader
      2 personalomsättning
    439 personen
     88 personens
    699 personer
     14 personerna
      2 personernas
      6 personers
      1 personhygienen
      1 personifierad
      1 personlift
     19 personlig
     31 personliga
      3 personligen
     19 personlighet
     18 personligheten
      2 personlighetens
      4 personligheter
      1 personlighetsavvikelser
      1 personlighetsdefekter
      9 personlighetsdrag
      1 personlighetsdraget
      1 personlighetsförändrade
      4 personlighetsförändring
      7 personlighetsförändringar
      1 personlighetsgenetik
      1 personlighetsgenetiken
      1 personlighetsgenetikens
      1 personlighetspsykologi
     58 personlighetsstörning
     24 personlighetsstörningar
      7 personlighetsstörningarna
      2 personlighetsstörningen
      1 personlighetsteori
      1 personlighetstyp
      1 personlighetstypen
      4 personlighetsutvecklingen
      1 personlighetsuveckling
     11 personligt
      1 personlyft
      1 personobj
     33 persons
      1 personsaneringsmedel
      1 personskada
      1 personskydd
      1 personskydds
      1 personuppgifter
     30 perspektiv
      1 perspektivenbr
      7 perspektivet
      1 perspektivtagande
      1 perspex
      1 perspiration
      1 persulcatus]
      1 pertaktin
      3 pertenue
      2 pertja
      5 pertussis
      1 pertussisgift
      1 pertussistoxin
      1 peruanska
      1 peruker
      1 perutz
      1 perversa
      1 perversion
      3 pes
      1 pescetarianism
      5 pessar
      1 pessargel
      5 pessimism
      1 pessimist
      1 pessimister
      2 pessimistisk
      1 pessism
     24 pest
      1 pestbakterie
      2 pestbakterien
      2 pestbakterier
      1 pestdoktor
      1 pestdoktorer
     53 pesten
      2 pestens
      1 pestepidemi
      1 pestepidemien
      1 pesticid
      1 pesticider
      1 pestilens
      5 pestis
      1 pestläkardräkt
      2 pestläkare
      1 pestlik
      1 pestloppan
      1 pestseptikemi
      1 pestsjukhus
      1 pestskråp
      1 pestsmittade
      1 pestutbrott
      1 pestvåg
      1 pestvatten
      3 pet
      5 peta
      1 petade
      2 petar
      1 petas
      1 petechier
      1 petekialt
      2 petekier
      8 peter
      1 petiolare
      1 petit
      1 petitmal
      1 petitmalepilepsi
      1 petning
      1 petrii
      1 petroleum
      1 petroleumprodukt
      1 petrovitj
      2 petscanning
      1 pettekniken
      1 petter
      2 pettersson
      2 peva
      2 peyronies
      1 pf
      2 pfenylendiamin
     27 pfizer
      4 pfizers
      1 pfk
      1 pg
     37 pga
      2 pglukos
      1 pglukosvärde
      2 pglukosvärdet
     38 ph
      1 phagein
      1 phagocytophilum
      1 phaléns
      1 phalloides
      1 phalloidin
      2 pharma
      1 pharmaceutical
      1 pharmaceuticals
      2 pharmacia
      1 pharmaciaprodukter
      1 pharmacop�a
      1 pharmacopœa
      2 pharmacopoeia
      1 pharmacopoeja
      1 pharmacy
      1 pharmakon
      3 pharynx
      1 phase
      1 phaselitanus
      1 phaseout
      1 phbalansen
      1 phberoende
      1 phbeteckning
      1 phd
      1 phellinus
      1 pherein
      1 phg
      1 phi
      1 phil
      4 philadelphia
      1 philadelphiakromosom
      1 philadelphiakromosomen
      1 philia
      5 philip
      1 philipp
      3 philippe
      1 philippine
     31 philips
      1 philishave
      1 philishaven
      2 philosophy
      4 phimosis
      1 phindikator
      1 phlebotomus
      1 phnivåer
      1 phnivåerna
      1 phnivån
      3 phobia
      2 phobos
      1 phocine
      1 pholiota
      1 phoma
      1 phoneutria
      1 phosphoenergon
      1 phreaking
      1 phrenicus
      2 phr�n
      1 phs
      3 pht
      1 phthiraptera
      1 phthisica
      2 phthisis
      1 phtls
      1 phtvålar
      1 phtvlphpv
     15 phvärde
      1 phvärden
      7 phvärdet
      1 phylicia
      1 physalia
      1 physalis
      2 physical
      2 physics
      4 physio
      2 phytolacca
      1 phytophthora
      2 pi
      1 pia
      1 pianisten
      1 piano
      1 pianosonat
      1 picasso
      1 picking
      1 picknick
      1 pickwick
      1 picoampere
      1 picornaviridae
      1 picornavirus
      1 picornavirusfamiljen
      1 pictogram
      1 picture
      1 pid
      1 piebaldism
      6 pierca
      2 piercad
      5 piercade
      1 piercades
      1 piercar
      1 piercare
      1 piercat
     11 piercing
      9 piercingar
      1 piercingarna
     10 piercingen
      5 pierre
      1 piezoelektrisk
      2 pigg
      1 pigga
      2 piggare
      2 piggen
      9 pigment
      4 pigmentceller
      1 pigmentcellerna
      1 pigmentcellstransplantationer
      2 pigmenten
      1 pigmenterade
      7 pigmentering
      1 pigmenteringen
      5 pigmentet
      2 pigmentförändring
      2 pigmentförändringar
      1 pigmentförluster
      1 pigmentlösa
      1 pigmentosa
      2 pigmentrubbningar
      1 pigtailkateter
      1 pikaktsignaleringsvägen
      1 piktogram
      4 pil
      1 pilar
      3 pilarna
      3 pilbågar
      1 pilbågen
      1 pilc
      1 pilegaard
      1 pilen
      1 pilgift
      1 pilgrimsfalk
      1 pilgrimsresor
      8 pili
      1 piliuttryck
      1 pilla
      1 pillar
     11 piller
      1 pillertrillande
      2 pillren
      1 piloerektion
      1 pilonidalcysta
      1 pilonidalsinus
      1 pilos
      1 pilot
      1 piloten
      2 piloter
      1 pilotglasögon
      1 pilotglasögonen
      1 pilotstudie
      1 pilprojektiler
      3 pilspets
      1 pilt
      1 pilus
      1 pimpinella
      1 pimpsten
      1 pinard
      1 piñata
      2 pincené
      1 pincenez
      7 pincett
      1 pincetten
      1 pincetter
      1 pineale
      1 pinealecysta
      3 pinel
      1 pingala
      1 pingviner
      1 pinjenötter
      2 pink
      1 pinka
      1 pinnar
      2 pinne
      1 pinocytos
      2 pinsamt
      3 pinta
      1 pinwale
      2 pinyin
      4 pionjär
      1 pionjärarbetet
      6 pionjärer
      2 pionjärerna
      1 pionjärinsatser
      1 pip
      7 pipa
      4 pipan
      5 pipande
      2 pipe
      1 piperidinderivat
      1 pipes
      1 pipig
      1 pipigt
     13 pipor
      1 piporna
      1 piprankeväxter
      1 piprensare
      1 piprökande
      2 piprökning
      1 pipstoppare
      1 piratkopiering
      1 piroxikam
      1 pirquet
      1 pirrande
      1 pirrningar
      1 pisiformis
      1 piska
      1 piskade
      1 piskades
      2 piskas
      1 piskmask
      1 piskor
      1 pisksnärt
      1 pisksnärtskador
      1 pisksnärtsskada
      1 pisksnärtsskador
      1 piso
      1 pissa
      1 pistaschnötter
      4 pistill
      1 pistillen
      1 pistiller
      3 pistol
      2 pitand
      2 pitands
      1 piteå
      1 piteälvarnas
      1 pitepaltar
      1 pitt
      1 pittha
      2 pittingödem
      1 pittoresk
      1 pittoreskt
      1 pituitary
      1 pityriasis
      1 pityrodeseksem
      2 pityrosporon
      1 pivmecillinam
      1 pixel
      1 pixie
      1 pixiebob
      1 pixlar
      1 pizza
      2 pjäs
      2 pka
      2 pkavärde
      1 pkryptorna
      5 pku
      1 pkudieten
      1 pkudrabbade
      1 pkutestet
      2 pl
     13 placebo
     10 placeboeffekten
      2 placeboeffekter
      1 placebogruppen
      1 placebokontrollerade
      1 placebopiller
      1 placebopreparat
      1 placeboresultaten
      1 placement
      2 placenta
      1 placentala
     11 placera
      8 placerad
     14 placerade
      6 placerades
     12 placerar
     58 placeras
      2 placerat
      3 placerats
     17 placering
      5 placeringen
      1 places
      1 placetett
     27 plack
      3 plackbildning
      1 placken
      1 plackens
      2 placket
      1 plackinnehåll
      1 plackmängden
      1 plackminskande
      2 plåga
      1 plågade
      2 plågades
      2 plågas
      1 plågat
      2 plågats
     14 plagg
      1 plaggen
      1 plagiat
      1 plagiatkontroll
      2 plågsam
      4 plågsamma
      2 plågsamt
      2 plague
     19 plan
      2 plana
      1 planare
      1 planchett
      2 plancks
      1 planen
      2 planer
      9 planera
      8 planerad
      8 planerade
      1 planerades
      1 planeraorganisera
      6 planerar
      3 planeras
      2 planerat
     13 planering
      5 planeringen
      1 planerings
      1 planeringsarbete
      5 planet
      1 plånet
      1 planlagd
      1 planlägga
      1 planläggning
      1 planlöst
      1 planmässigt
      1 planschetten
      1 plant
      3 planta
      1 plantager
      5 plantan
      1 plantans
      1 plantar
      1 plantarfascia
      1 plantarfascian
      2 plantarfasciasenan
      7 plantarfasciit
      1 planten
      1 plantera
      1 planteras
      1 plantering
      2 planteringar
      1 planteringstid
      7 plantor
      2 plantorna
      1 plantz
      1 plaques
     20 plasma
      1 plasmacell
      3 plasmaceller
      2 plasmacellerna
      1 plasmacellsmyelom
      1 plasmaelektrofores
      1 plasmaersättningsmedel
      1 plasmaferes
      1 plasmakomponenter
      1 plasmakoncentration
      1 plasmakoncentrationen
      1 plasmakoncentrationer
      1 plasmakoncentrationerna
      1 plasmalemma
      2 plasmamembran
      5 plasmamembranet
      1 plasmamembranets
      5 plasman
      1 plasmanivåer
      1 plasmapelare
      6 plasmaproteiner
      1 plasmaproteinerna
      1 plasmaproteinet
      1 plasmaproteinfraktionering
      1 plasmavolym
      2 plasmid
      3 plasmidburen
      1 plasmidburna
      2 plasmider
      1 plasmiderna
      1 plasmidmedierad
      3 plasmin
      2 plasminogen
      1 plasminogenaktivator
      1 plasmodier
      2 plasmodiophora
      1 plasmodiophoromycota
      1 plasmodium
      1 plasmodiumsläktet
      1 plassein
     30 plast
      1 plastade
      1 plastbågar
      2 plastbehållare
      1 plastbygel
      1 plastbyxor
      1 plastdetaljer
     11 plaster
     22 plåster
      2 plasterna
      1 plastförpackningen
      1 plastfyllning
      2 plastglas
      1 plastglaset
      1 plastgruppen
      1 plastgummi
      4 plasticitet
      1 plasticiteten
      2 plastik
      1 plastikirurgin
      1 plastikkirgiskt
      2 plastikkirurg
      2 plastikkirurgen
      1 plastikkirurger
     18 plastikkirurgi
      5 plastikkirurgin
      6 plastikkirurgisk
      1 plastikkirurgiska
      1 plastikkirurgiskt
      1 plastikoperationer
      1 plastikopereration
      1 plastikos
      3 plastisk
      1 plastiska
      1 plastiskt
      1 plastkatetrar
      1 plastklädnypor
      1 plastkondomer
      1 plastkoppar
      1 plastkroppar
      2 plastmaterial
      1 plastmattor
      1 plastmöbler
      1 plastpåsar
      1 plastpåsarnas
      2 plastpåse
      1 plastremsa
      3 plåstret
      2 plastringar
      1 plaströr
      1 plastrum
      1 plastscintillatorer
      1 plastsida
      1 plastskaft
      1 plastskal
      1 plastskålar
      1 plastskena
      1 plastslang
      1 plastsula
      1 plasttallrikar
      1 plasttuben
      1 plåta
      1 platanthera
      1 plåtbitar
      1 plateau
      1 platelet
      5 platon
      1 platoniska
      1 platonismen
      1 platons
      1 plåtränna
     93 plats
      1 platsanalys
      1 platsbrist
     18 platsen
      1 platsens
     66 platser
      2 platserna
      1 platsproblem
      1 platsteorin
     10 platt
     14 platta
      1 plattade
      1 plattan
      2 plattar
      2 plattare
      3 plattas
      2 plattepitel
      2 plattform
      1 plattformen
      2 plattfot
      1 plattfota
      1 plattfotheten
      2 plattmaskar
      1 plattmaskarna
     13 plattor
      2 plattparet
      1 platytaenium
      1 plavix
      2 plc
      2 pleconaril
      1 plecostachys
      1 plectranthus
      1 plenipotentiär
      1 pleokroism
      1 pletysmograf
      4 pleura
      1 pleuracancer
      1 pleurahålan
      1 pleural
      4 pleuran
      3 pleuraplack
      1 pleuraplacken
      1 pleuratappning
      1 pleuratrycket
      2 pleurautgjutning
      1 pleurautgjutningar
      1 pleuravätska
      1 pleuritisk
      1 pleuritiska
      1 pleuropulmonära
      4 plexiglas
      4 plexus
      1 p�li
      1 pliktverket
      2 plinius
      1 pljudet
      9 plocka
      1 plockad
      1 plockades
      2 plockar
      7 plockas
      3 plockning
      1 ploetz
      1 plommon
      1 plotinos
      1 plötligt
     28 plötslig
      5 plötsliga
      1 plötsligen
     43 plötsligt
      1 plotta
      1 plottar
      1 plottas
      4 plugg
      1 plugga
      1 pluggarna
      1 pluggskivling
      1 plumbsticks
      1 plumbum
      4 plur
      6 plural
      1 pluralis
      7 plus
      1 plusgrader
      1 pluspol
     24 plutonium
      1 plutoniumisotoper
     14 plutoniums
      1 plymer
      1 plymouths
      2 pm
      1 pmitrale
      4 pmma
      4 pms
      1 pmsbesvär
     13 pmt
      1 pmtbehandlingsmetod
      1 pmtmetod
      1 pmtmetoden
      1 pmtmetoder
      1 pmtutbildning
      1 pnets
      1 pneumatologer
      1 pneumatologi
      3 pneumatologin
      1 pneumatologiska
      2 pneumocystis
      1 pneumocystispneumoni
      1 pneumocyternas
      1 pneumokocken
      1 pneumokockens
     23 pneumokocker
      2 pneumokockerna
      4 pneumokockinfektioner
      1 pneumokockkonjugatvaccin
      3 pneumokockmeningit
      2 pneumokockpneumoni
      1 pneumokockpolysackaridvaccinet
      1 pneumokocksjukdom
      3 pneumokockvaccin
      2 pneumokonios
      1 pneumonektomi
     31 pneumoni
      3 pneumonia
     15 pneumoniae
      1 pneumonifynden
      1 pneumonii
      1 pneumonin
      4 pneumonit
      6 pneumophila
      3 pneumothorax
     11 po
     18 poäng
      1 poängbedömining
      5 poängen
      1 poänglösa
      1 poängresultatet
      1 poängsätta
      1 poängsätter
      1 poängskalor
      1 poängsmoment
      1 poängsumma
      1 poängsumman
      1 poängsystemet
      1 poängtal
      1 poängtera
      1 poängterade
      3 poängterar
      1 pocker
      4 podiatri
      1 podiatric
      4 podiatriker
      1 podiatrikerna
      1 podiatrin
      1 podiatry
      1 podoconiosis
      1 podocytisus
      1 podofyllotoxin
      1 poecilia
      1 poem
      3 poesi
      1 poesins
      4 poeten
      2 poetiska
      1 poetry
      1 pofloden
      2 pogosta
      2 pogostasjuka
      1 poiein
      1 point
      1 points
      5 poison
     65 pojkar
      2 pojkarmän
     12 pojkarna
      1 pojkarnas
      2 pojkars
     16 pojke
     16 pojken
      4 pojkens
      1 pojkfoster
      1 pojkfostrets
      1 pojkgiftermålen
      1 pojkmetoder
      1 pojkvänner
      1 poker
      1 pokermaskiner
      1 pöl
      1 pölar
      2 polär
      3 polära
      1 polarisation
      1 polarisationsfilter
      2 polariserade
      1 polaritet
      1 polaroidsolglasögon
      1 polarregioner
      2 polarregionerna
      1 polärt
      1 póleis
     15 polen
      1 poler
      1 polerar
      3 poleras
      4 police
      5 policy
      1 policydokument
      4 policyn
      1 poliklinikpatienter
      1 poliklinisk
      1 polikliniskt
      3 polio
     20 polis
      1 pólis
      1 polisanmäldes
      1 polisarbete
      1 polisbåtar
      2 polisbilar
      1 polisbricka
      1 polisdistrikt
      1 polisdistriktet
     38 polisen
      6 polisens
      5 poliser
      2 polisers
      1 polisfordon
      1 polishästar
      1 polishelikoptrar
      1 polisiär
      6 polisiära
      1 polisingripande
      1 polisinsatser
      2 poliskår
      7 poliskårer
      1 poliskårerna
      1 poliskommissarie
      1 poliskonstapel
      1 poliskunder
      1 polislegitimation
      1 polislegitimationen
      1 polismakt
      1 polisman
      1 polismannen
      1 polismästare
      1 polismotorcyklar
      2 polismyndigheten
      1 polismyndigheterna
      1 polisorgan
      1 polisradio
      1 polisstaten
      1 polisstationer
      1 polisstyrka
      1 polisstyrkan
      1 polisuniform
      1 polisväsen
      1 polisväsenden
      3 polisväsendet
      1 politeia
      1 politia
      7 politik
      1 politiká
      3 politiken
      8 politiker
      3 politikern
      1 politikområdet
      1 politikós
      7 politisk
     20 politiska
      1 politiske
      7 politiskt
      1 polkärnorna
      2 polkropp
      1 polkroppar
     26 pollen
      1 pollenallergen
      1 pollenallergenet
     10 pollenallergi
      3 pollenallergiker
      1 pollenanalys
      1 pollenet
      2 pollenkorn
      3 pollenkornen
      1 pollenkornens
      2 pollenkornet
      1 pollenmediciner
      1 pollensäsong
      1 pollensäsongen
      1 pollenslang
      2 pollenslangen
      1 pollenslangscell
      1 pollinatörer
      1 pollineras
      5 pollinering
      1 pollineringen
      2 pollution
      1 pollutioner
      1 polo
      7 polonium
      1 poloniumisotoper
      1 poloniumisotoperna
      1 polske
      1 polus
      2 poly
      1 polycykliskt
      1 polycystisk
      1 polycystiska
      7 polycystiskt
      1 polycytemi
      2 polydaktyla
     10 polydaktyli
      2 polydaktylin
     12 polydipsi
      1 polyelektrolyter
      1 polyembryoni
      3 polyester
      1 polyfenoler
      1 polyfenylenoxid
      2 polyfyletiska
      1 polygama
      1 polygenetisk
      1 polyglutaminkedja
      1 polyglutaminkedjan
      1 polyglykolsyra
      1 polygrafisk
      1 polyhydroxylerat
      1 polykarbonat
      2 polyklorerade
      1 polyklorering
      2 polykromatisk
      2 polymer
      1 polymerase
      5 polymeraskedjereaktion
      1 polymeren
      4 polymerer
      1 polymerfibrer
      1 polymerform
      1 polymeriseras
      1 polymerisering
      1 polymermaterial
      1 polymernätverket
      1 polymethylmethacrylatebågar
      1 polymetylmetakrylat
      4 polymorfa
      2 polymorfismer
      1 polymorphus
      6 polymyosit
      1 polymyxin
      1 polynesien
      1 polynesier
      1 polynesiska
      2 polyneuropati
      5 polyp
      3 polypen
      1 polypens
      3 polypeptid
      5 polypeptider
      1 polypeptidernas
      2 polypeptidhormon
      1 polypeptidkedja
      1 polypeptidkedjor
     16 polyper
      1 polyphyllus
      1 polyporales
      1 polypropylen
      1 polyq
      1 polyqkedjan
      4 polysackarid
      1 polysackariddel
      1 polysackariddelen
      2 polysackariden
      3 polysackarider
      1 polysackariderna
      2 polysackaridkedjorna
      3 polysomnografi
      2 polysomnografier
      1 polysorbat
      3 polyspermi
      1 polystyren
      1 polystyrensulfonat
      1 polyteistiska
      1 polyuretan
     16 polyuri
      1 polyuria
      3 polyurin
      1 polyvinylklorid
      1 pombe
      8 pomc
      1 pomcbrist
      1 pomcgenen
      1 pomcnullsyndromet
      2 pomcs
      2 pompejus
      1 ponds
      1 ponoconiosis
      5 pons
      1 ponseti
      1 ponsetimetoden
      1 ponsvinkeltumör
      2 ponti
      1 pontiac
      2 pontiacfeber
      2 pontos
      1 pontsaintesprit
      1 poolen
      2 pop
      1 popgruppen
      1 poppel
      1 poppelsläktet
      2 popper
      1 poppers
     24 populär
     18 populära
      1 populärare
      2 populärast
      3 populäraste
      2 populariserade
      3 populariserades
      9 popularitet
      1 popularitetsskäl
      6 populärkultur
      5 populärkulturen
      3 populärnamn
     30 populärt
      1 populärvetenskapligt
     22 population
     18 populationen
      1 populationens
      9 populationer
      1 populationsgenetik
      1 populationsstudier
      1 populationstrenden
      1 populous
      1 por
      1 porath
      1 porbitalerna
      8 porer
      2 porerna
      1 porfobilinogen
      7 porfyri
      4 porfyrier
      3 porfyrierna
      2 porfyrin
      1 porfyrindelar
      3 porfyriner
      1 porfyrinerna
      3 porfyrinet
      1 porinproteinerna
      1 porinproteinet
      1 pormaskar
      1 pörn
      1 pornografi
      1 pornografiberoende
      2 poröst
      1 porphyra
      1 porro
      1 porros
      1 porrstjärnor
      1 pors
      2 porslin
      1 porslinsguden
      1 porslinssked
      2 porslinsskrammel
      1 porsystemens
      2 port
      3 porta
      2 portabel
      1 portådern
      1 portådersystem
      1 portae
      2 portahypertension
      1 portakretslopp
      1 portakretsloppet
      4 portal
      1 portalfigur
      1 portalhypertoni
      1 portalområderna
      2 portar
      1 portasystem
      2 portasystemet
      1 portasystemisk
      1 portavenen
      1 pörte
      1 portefaix
      4 portfölj
      2 portföljen
      1 portioner
      1 portionera
      1 portionerar
      1 portionsförpackad
      4 porträtt
      1 porträtten
      1 porträtteras
      1 porträttkonst
     19 portugal
      1 portugaltyskland
      1 portugis
      1 portugiser
      2 portugisisk
      3 portugisiska
      1 portugisiske
      1 portvakt
      5 portvenen
      1 portvinsfärgad
      1 portvinstå
      1 poser
      3 pösiga
     19 position
      3 positionen
      6 positioner
      1 positionerade
      1 positioneringen
      4 positionerna
      1 positioning
      1 positionsangivelse
      1 positionsberoende
     58 positiv
     82 positiva
      8 positive
     40 positivt
      3 positron
      1 positronemissionstomografi
      1 positronemissiontomografi
      1 positronen
      1 positroner
      1 possehl
      2 post
      1 posten
      2 postencefalitiskt
      2 poster
      3 posteriora
      1 posteriori
      1 posteriort
      1 postexponeringsbehandling
      2 postexpositionsprofylaktisk
      1 postexpositionsprofylax
      1 postgangliona
      1 postgymnasial
      1 posthallucinatorisk
      1 posthepatisk
      2 postherpetisk
      1 posthypnotisk
      2 postinfektiös
      1 postlunchdip
      1 postmenopaus
      1 postmenopausala
      1 postnataldepressioner
      2 postoperativa
      1 postoperativt
      1 postorder
      1 postpartum
     13 postpartumdepression
      5 postpartumdepressioner
     11 postpartumpsykos
      4 postpartumpsykoser
      1 postpartumtyreoidit
      1 postpeak
      1 postpunk
      1 postrema
      2 postschizofren
      1 postspinal
      1 postsynaps
      1 postsynapsens
      2 postsynaptisk
      7 postsynaptiska
      8 posttraumatisk
     13 posttraumatiskt
      1 postulerar
      1 postum
     12 potatis
      1 potatisåkrar
      2 potatisbladmögel
      1 potatischips
      1 potatissläktet
      1 potatisväxt
      6 potatisväxter
      5 potens
      3 potensen
      2 potenser
      1 potensproblem
      6 potent
      3 potenta
      1 potentare
      1 potentaste
      7 potential
      1 potentialen
      1 potentialminimum
      1 potentialskillnaden
      2 potentiell
     10 potentiella
     28 potentiellt
      1 potentiera
      1 potentierade
      1 potentiering
      1 potentieringar
      1 potientellt
      1 potomani
      4 potta
      1 potter
      1 potts
      2 pouch
      1 pourprejpgfullvuxna
      1 pousette
      1 pousettes
      1 povel
      1 povidonjod
      1 pow
      1 poweryoga
      1 pox
      1 poxviridae
      2 poxvirus
      1 pozzed
      1 ppd
      1 ppg
      1 ppi
     23 ppiller
      1 ppilleranvändning
      1 ppillerbehandlingen
      2 pplåster
      6 ppm
      1 ppmdirekt
      1 ppo
      1 pprotrombinkomplex
      1 ppulmonale
      2 pqtid
      1 pra
      1 pr�a
      1 practice
      1 practitioner
      3 praecox
      1 praetoria
      2 praetoriangardet
      1 praevalens
      1 praevia
      1 prag
      2 prägel
      3 prägla
      4 präglad
      8 präglade
      2 präglades
      3 präglar
     13 präglas
      1 präglats
      1 pragmatik
      2 pragmatiska
      1 pragmatiskt
      1 pragmatism
      1 prakiskt
      1 praktfull
      2 praktfulla
     15 praktik
     36 praktiken
      2 praktiker
      1 praktikerna
      1 praktikterminen
      1 praktikterminerna
      1 praktisera
      1 praktiserad
      2 praktiserades
      3 praktiserande
      1 praktiserar
      5 praktiseras
      1 praktiserat
     12 praktisk
     19 praktiska
      1 praktiskakliniska
     29 praktiskt
      1 praktos
      3 prana
      1 pranan
      3 pranayama
      1 präriehundar
      1 prärievarg
      1 prärievargar
      2 präst
      1 prästämbete
      3 prästen
      6 präster
      1 prästerna
      1 prästerskapet
      1 prästerskapets
      1 prästliknande
      1 prästnäsduk
      1 prästs
      5 prat
     15 prata
      2 pratade
     13 pratar
      1 pratat
      1 pravachol
      1 praxinoskopet
     10 praxis
      2 praziquantel
      1 prazol
      3 pre
      1 prebiotika
     60 precis
      2 precisera
      1 preciserade
     11 precision
      2 precisionen
      1 precisionsdiagnostisk
      1 precisionsinstrument
      1 precisionsmätningar
      1 precisionsstrålningsteknik
      1 precolumbian
      1 precolumbianska
      1 precordiala
      1 precox
      1 predatorer
      1 predestinera
      1 predicera
      1 predikningar
      2 prediktionsregler
      1 prediktiva
      1 prediktorerna
      3 predisponerad
      2 predisponerade
      5 predisposition
      1 predispositioner
      1 prednisolon
      3 predominantly
      8 preeklampsi
      1 preembryoperioden
      2 preexcitation
      1 preexcitationen
      2 preferens
      2 preferenser
      1 preferenserna
      6 prefix
      2 prefixet
      4 prefrontala
      1 prefrontalcortex
      1 prefrontalloberna
      1 pregabalin
      1 pregnancy
      2 pregnenolon
      1 prehallux
      1 prehepatisk
      2 prehospital
      1 prehospitalt
      2 preimplantatorisk
      1 prejudicerande
      1 prekapillära
      3 prekursor
      2 prelamin
      2 preliminär
      3 preliminära
      1 preload
      2 preludin
      4 prematur
      6 prematura
      1 prematurfödelse
      1 prematurity
      2 premenopausal
      4 premenstruell
      1 premenstruella
      3 premenstruellt
      1 premierna
      1 premisser
      1 premiumprodukter
      1 premotoriska
      1 prenumererad
      1 preoperativa
     81 preparat
     13 preparaten
     35 preparatet
      2 preparatets
      1 preparatgrupp
      2 preparation
      1 preparationer
      2 preparativ
      1 preparats
      1 preparera
      2 preparerade
      1 prepareras
      1 preparerat
      1 prepatellarbursit
      1 preposition
      1 preprohypokretin
      1 preproinsulin
      1 preproinsulinet
      5 prepsykos
      3 prepsykosen
      2 prepsykosens
      3 prepsykoser
      1 prepsykotiska
      1 prepubertala
      1 prepuberteten
      1 presbyoper
      5 presbyopi
      1 presenil
      1 presenningar
      1 presens
      1 present
      6 presentation
      1 presentationen
      1 presentations
      6 presentera
      1 presenterad
      6 presenterade
      4 presenterades
      9 presenterar
      7 presenteras
      1 presenterat
      5 presenterats
      1 president
      5 press
      4 pressa
      3 pressade
      1 pressades
      8 pressar
     18 pressas
      3 pressat
      1 pressduk
      1 pressen
      1 pressetiska
      1 pressgjutas
      1 pressjärn
      2 pressjärnet
      1 pressmeddelande
      1 pressning
      7 pressure
      6 prestanda
      1 prestandaförmågan
      7 prestation
      4 prestationen
      1 prestationer
      1 prestationerna
      2 prestationsångest
      3 prestationsförmåga
      2 prestationsförmågan
      1 prestationsmotivation
      2 prestera
      8 presterade
      1 presterande
      1 presterar
      1 presterat
      1 prestigefulla
      1 prestigefyllda
      1 presynaps
      2 presynapsen
      3 presynaptisk
      4 presynaptiska
      3 pretibialt
      2 preussen
      1 preussens
     18 prevalens
     16 prevalensen
      1 prevalensuppskattning
      1 prevalensuppskattningar
     25 prevention
      1 preventionref
      2 preventionsmetod
      2 preventiv
      4 preventiva
      1 preventive
     34 preventivmedel
      1 preventivmedels
      1 preventivmedelsbehov
      1 preventivmedelsmottagning
      1 preventivmedelsrådgivning
      3 preventivmedlen
      2 preventivmedlet
      3 preventivmetod
      2 preventivmetoden
      2 preventivmetoder
      4 preventivt
      1 preventol
      1 prév�ts
      1 priapi
     22 priapism
      2 priapos
      2 prick
      1 pricka
     12 prickar
      1 prickensåret
      1 prickig
      1 prickskyttegevär
      9 pricktest
      1 pricktesten
      2 pricktester
      3 priessnitz
      1 priest
      1 priestley
      2 primal
      1 primalakulär
      1 primalinstitutet
      1 primalskriket
      2 primalterapi
      3 primalterapin
      1 primalterapins
     50 primär
     45 primära
      1 primärfallet
      2 primärgranula
      1 primärinfektion
      1 primärkällan
      1 primärkänsla
      1 primärläkare
      1 primärspole
     27 primärt
      1 primärtumör
      1 primärtumören
      1 primärtumörer
      2 primärvård
      7 primärvården
      1 primary
      1 primatarter
     13 primater
      4 primitiva
      1 primitivare
      1 primitivaste
      2 primitivism
      2 primitivt
      1 primolut
      1 primroten
      1 primum
      1 princeton
     38 princip
     20 principen
     21 principer
      5 principerna
      1 principiell
      2 principiella
      2 principiellt
      1 principle
      4 pring
      2 pringar
      1 pringarna
      1 pringen
      1 prins
      1 prinsessan
      1 prinskorv
      1 prinskorvsliknande
      1 print
      1 printerval
      4 prion
     11 prioner
      3 prionerna
      1 prionet
      1 prionprotein
      2 prionsjukdom
      1 prionsjukdomar
      3 prionsjukdomarna
      1 prionsjukdomen
      1 priori
      1 prioritera
      4 prioriterar
      6 prioriteras
      2 prioriterat
      3 prioritering
      2 prioriteringar
      1 prioritet
      9 pris
      1 prisade
      1 prisades
      3 prisbild
      5 priser
      2 priserna
     14 priset
      1 prisklasserna
      1 prislappar
      3 prisma
      1 prispengarna
      1 prissättningsstrategier
      1 pristagare
      1 prithvi
     15 privat
     23 privata
      1 privathem
      1 privatimport
      2 privatkök
      1 privatkunder
      1 privatperson
      1 privatpersonen
      7 privatpersoner
      1 privatskolaför
      1 privattandläkare
      1 privilegiebrev
      1 privilegiehandel
      1 privilegiet
      2 privilegium
     10 pro
      1 proactiv
      1 proactive
      7 proana
      1 proanasajter
      2 prob
      1 probably
      1 proben
      1 prober
     24 probiotika
      1 probiotikabakterier
      1 probiotikabakterierna
      1 probiotikaforskningen
      6 probiotikan
      2 probiotikans
      1 probiotikapiller
      1 probiotikor
      2 probiotisk
      5 probiotiska
    338 problem
      1 problemartat
      1 problemataxxxi
     13 problematik
      7 problematiken
      1 problematiseras
      8 problematisk
      9 problematiska
      7 problematiskt
      3 problembeteenden
      1 problembeteendena
      1 problembilden
     31 problemen
     42 problemet
      1 problemfria
      1 problemkonsumenter
      1 problemläkemedlet
      3 problemlösning
      1 problemlösningsförmågor
      1 problemmedvetenhet
      1 problemområdet
      2 problems
      1 problemstörningar
      1 probnp
      1 probnukleinsyrekedjor
      1 procedirer
      7 procedur
      8 proceduren
      1 procedurer
      1 proceedings
    204 procent
      5 �procent
      1 procentantalet
      4 procenten
      3 procentenheter
      2 procenthalt
      2 procentig
      4 procents
      2 procentsats
      1 procenttal
      2 procenttalet
      1 procentuella
      1 procentvärde
      1 procera
     95 process
      1 processandet
      2 processas
     52 processen
     39 processer
      1 processerad
      3 processerna
      1 processfärdigheterna
      1 processing
      1 processvärme
      1 procter
      1 proctor
      1 prodentis
      1 prodesse
      8 prodrom
      1 prodromalstadium
      1 prodromen
      1 prodromsymtomen
      1 prodrug
      1 prodrugs
      4 producenter
     57 producera
      4 producerad
     10 producerade
      5 producerades
     93 producerar
     57 produceras
      3 producerat
      6 producerats
      1 product
      3 products
      1 produker
     21 produkt
     18 produkten
      4 produktens
     91 produkter
     12 produkterna
      1 produkters
      1 produktervaror
      1 produktgodkännande
      1 produktgrupper
     57 produktion
     43 produktionen
      1 produktionsbortfall
      1 produktionsdjur
      1 produktionslinjer
      1 produktionsmetoder
      1 produktionsnivåerna
      1 produktionsomgång
      1 produktionssorterna
      1 produktionstekniken
      3 produktiv
      1 produktivitet
      1 produktkontroll
      1 produktkontrollen
      1 produktnamnet
      1 produktresumé
      1 produktspecifik
      1 produktutvecklingspartnerskap
      1 proenzym
      3 prof
      1 profana
      1 professing
      3 profession
      1 professionalisering
      8 professionell
      8 professionella
      5 professionellt
      1 professioner
     27 professor
      1 professorer
      1 professorerna
      4 professorn
      1 professur
      1 professuren
      2 professurer
      1 professurerna
      1 profeten
      1 profeternas
      1 profetior
      2 proffs
      1 proffsdansare
      5 profil
      1 profile
      3 profiler
      1 profilområde
      1 profunda
      1 profylaktik
      6 profylaktisk
      2 profylaktiska
      2 profylaktiskt
      3 profylax
      1 progenitor
      3 progenitorcell
      2 progenitorceller
      9 progeri
      6 progeria
      1 progerin
      1 progerisjuka
      1 progerisjukas
      1 progerisyndromen
      1 progestagen
     29 progesteron
      1 progesteronet
      1 progesteronfasen
      1 progesteronhalten
      1 progesteronhämmare
      1 progesteronpreparat
      1 progesteronreceptorer
      1 progesteronvärden
      1 progeston
     40 prognos
     37 prognosen
      1 prognoserna
      1 prognostisera
      1 prognostisk
      2 prognostiskt
     30 program
      1 programkod
      4 programme
      4 programmen
      1 programmens
      1 programmera
      3 programmerad
      1 programmerade
      1 programmeras
      1 programmerat
     13 programmet
      1 programmets
      6 programvara
      1 programvaran
      1 progredierande
      1 progredierar
      1 progress
      4 progression
      1 progressionen
      6 progressiv
     14 progressiva
      3 progressivt
      5 prohibition
      1 prohibitionism
      1 prohibitionister
      1 prohibitionisters
      1 prohibitionistiskt
      5 prohormon
      4 prohormoner
      1 prohormonkonvertaser
      3 proinflammatoriska
      3 proinsulin
      3 proinsulinet
      2 projection
      9 projekt
      1 projektarbeten
     12 projektet
      6 projektion
      5 projektioner
      1 projektionsavbildning
      1 projektionsmetod
      1 projektionsriktningen
      1 projicera
      1 projicerad
      1 projicerade
      1 projicerar
      1 projiceras
      2 projicering
      2 prokain
      1 prokalcitonin
      3 prokaryota
      1 prokaryoter
      1 proktolog
      1 proktologi
      1 proktoskop
     21 prolaktin
      1 prolaktinet
      1 prolaktinets
      1 prolaktinhämmande
      5 prolaktinnivåer
      1 prolaktinnivåerna
      2 prolaktinom
      1 prolaktinproduktionen
      1 prolaktinreceptorer
      1 prolamin
      1 prolaminet
      1 prolaps
      3 proliferation
      1 proliferativa
      1 prolin
      1 promenad
      4 promenader
      1 promenera
      1 promenerar
      2 promia
      3 promille
      1 promilles
      3 promiskuitet
      1 promoe
      1 promotades
      1 promotion
      1 promyelocyte
      4 pronation
      1 pronationens
      1 pronerar
      1 pronomroblasten
      1 pronormoblast
      1 proopiomelanokortin
      1 prop
      1 propagerade
      1 propan
      3 propanol
      5 propantriol
      2 propen
      1 propensulfensyra
      1 proper
      1 properties
      1 property
      1 propiomazin
      1 propionsyra
      4 propofol
      7 proportion
      1 proportional
      5 proportionell
      2 proportionellt
      4 proportioner
      2 proportionerna
      2 proposition
      9 propp
      3 proppar
      2 proppbildning
      1 proppbildningsrisk
      9 proppen
      2 propplösande
      1 proppmätte
      2 propria
      1 propylenglykol
      1 propylhexedrin
      1 propylpentansyra
      1 prosit
      9 prosopagnosi
      1 prosopon
      1 prospektering
      1 prospekteringsbolag
      2 prospektiv
      1 prósstata
      5 prostaglandiner
      1 prostaglandinhämmande
      1 prostaglandinhämmarna
      1 prostait
     20 prostata
     44 prostatacancer
      1 prostatacancerpatienter
      1 prostatafall
      1 prostataförstoring
      2 prostatahyperplasi
      1 prostatakörtel
      1 prostatakörteln
      1 prostatakörtelns
      1 prostatamassage
      7 prostatan
      1 prostatans
      1 prostataproblem
      3 prostatasekret
      1 prostatasekretet
      1 prostatasjukdomar
      4 prostataspecifikt
      3 prostatektomi
     10 prostatit
      1 prostatitdiagnoser
      1 prostituerad
      5 prostituerade
      6 prostitution
      2 protagonist
      1 protagonisten
      1 protagonistens
      1 protallier
      1 protaminer
      1 proteas
      2 proteaser
      2 protection
    108 protein
      1 proteinaggregat
      1 proteinämnen
      1 proteinansamlingar
      1 proteinberikad
      1 proteinbildningen
      1 proteinbrist
      1 proteindelen
      1 proteinen
     82 proteiner
      8 proteinerna
      1 proteinernas
      2 proteiners
     42 proteinet
      1 proteinets
      1 proteinfamiljen
      2 proteinfattig
      2 proteinfattiga
      2 proteinförgiftning
      2 proteinfragment
      4 proteinhalt
      3 proteinhalten
      1 proteinhormon
      3 proteininnehåll
      2 proteinintag
      1 proteinintaget
      2 proteinkapsel
      1 proteinkedjan
      2 proteinkedjor
      1 proteinklister
      2 proteinkomplex
      1 proteinkomplexen
      1 proteinkristaller
      1 proteinnedbrytning
      1 proteinnivåer
      1 proteinprodukt
      4 proteinrik
      2 proteinrika
      1 proteinrikt
      1 proteins
      1 proteinsammansättningar
      6 proteinsyntes
      6 proteinsyntesen
      1 proteintillskott
      1 proteintillverkning
      2 proteinuri
      1 proteinveckning
      1 proteobacteria
      1 proteobakterier
      2 �proteobakterierna
      1 proteoglycans
      1 proteoglykaner
      1 proteolys
      1 proteolysen
      1 proteolytiska
      3 proteolytiskt
      1 proteos
      9 protes
      5 protesen
      1 protesens
      8 proteser
      2 proteserna
      1 proteskirurgi
      1 protesoperation
      2 protest
      1 protestantiska
      3 protester
      1 protesterade
      1 protesterande
      1 protesthandling
      1 protestillverkare
      3 protetik
      1 protetiker
      1 protetiska
      2 proteus
      1 prothorax
      1 proto
      1 protoindoeuropeiska
      1 protoklorofyllid
      1 protokollavkodningar
      1 protokollet
      1 protokollförande
      1 protolyseras
      6 protoner
      1 protonerat
      1 protongradienten
      6 protonpumpshämmare
      2 protonpumpshämmarna
      1 protonterapi
      1 protoonkogen
      2 protoonkogenen
      2 protoonkogener
      1 protopic
      1 protoplasma
      1 protoporfyrin
      1 prototypen
      2 protozoa
      1 protozoen
      6 protozoer
      1 protozoisk
      1 protozooer
      4 protrombin
      1 proust
     38 prov
      5 prova
     10 pröva
      3 provade
      5 prövade
      2 prövades
      1 provar
      1 prövar
      1 prövaren
      2 provas
      9 prövas
      2 provat
      2 prövat
      2 provats
      6 prövats
      1 provdnat
     15 prover
      3 proverna
     20 provet
      1 provexcision
      2 provfiske
      1 provide
      1 providencekorsetten
      1 provins
      1 provinsamling
      4 provinsen
      1 provinser
      1 provinserna
      1 provinsialläkarväsendet
      1 provisional
      1 provisoriskt
      1 provisorsexamen
      1 provlämning
      1 provmaterial
      1 provmetoderna
      1 provning
     16 prövning
     11 prövningar
      2 prövningarna
      2 prövningen
      1 prövningsdata
      1 prövningsinstansen
      1 prövningstillstånd
      3 provocerad
      5 provocerade
      1 provocerande
      2 provocerar
      4 provokation
      2 provokationer
      1 provokativ
      4 provrör
      2 provrören
      1 provrörsbarn
      1 provsticka
      3 provsvar
      1 provsvaren
     17 provtagning
      1 provtagningar
      3 provtagningen
      1 provtagningsröret
      1 provtavlan
      1 prowazekii
      1 proximala
      1 proximalt
      3 prpc
      2 prpsc
      1 prunus
      1 pruritic
      1 prusa
      2 prusiner
      1 prustrot
      1 prutt
      1 pruttkudde
      1 pruttljud
      1 prydd
      1 prydda
      1 pryddes
      1 prydliga
      2 prydnad
      1 prydnader
      1 prydnadsbuske
      1 prydnadsföremål
      1 prydnadsspänne
      9 prydnadsväxt
      5 prydnadsväxter
      1 pryds
      1 pryglade
      1 pryglades
      1 pryl
      1 psa
      1 psaprovtagning
      2 pse
      1 psekret
      1 pseudoafaki
      2 pseudoakromegali
      1 pseudoanafylaxi
      1 pseudoartros
      1 pseudocapsicum
      1 pseudocicera
      1 pseudocoelomata
      1 pseudodemens
      1 pseudodyskalkyli
      1 pseudoefedrin
      2 pseudogikt
      1 pseudohallucination
      1 pseudohermafroditism
      1 pseudokrupp
      1 pseudolaglig
      6 pseudomonas
      2 pseudomorf
      1 pseudonaja
      1 pseudonarcissus
      1 pseudoneurologiska
      1 pseudonym
      1 pseudoord
      1 pseudoteorier
      1 pseudoterranova
      1 pseudotorticollis
      8 pseudovetenskap
      1 pseudovetenskaplig
      2 pseudovetenskapliga
      1 pseudovetenskapligt
      1 psg
      1 psilocybin
      3 psittaci
      1 psittacinafåglar
      1 psittacos
      1 psittakos
      1 psocoptera
      1 psoralea
      6 psoralen
      1 psoralener
     15 psoriasis
      1 psoriasisartit
      8 psoriasisartrit
      1 psoriasisbehandling
      1 pspruta
      1 psprutan
      3 pstav
      3 pstavar
      5 pstaven
      1 psv
      4 psvt
      1 psych�
      3 psyche
      1 psyché
      1 psychein
      3 psychiatric
      1 psychoanalysis
      1 psychoanalytical
      1 psychobiology
      1 psychological
      1 psychometric
      1 psychopathology
      1 psychopetem
      2 psychosis
      1 psychotherapy
      3 psykasteni
      1 psykasteniskarubbningar
     15 psyke
      1 psykedelisk
      4 psykedeliska
      1 psykedeliskt
     15 psyket
      1 psykhe
      1 psykiaktrisk
      7 psykiater
      1 psykiaterförbundet
      9 psykiatern
      1 psykiaterns
      2 psykiatrer
      2 psykiatrerna
     20 psykiatri
      1 psykiatrifältet
      6 psykiatriker
      4 psykiatrikern
      1 psykiatrikernas
      1 psykiatrikritik
      1 psykiatrikritiken
     30 psykiatrin
      7 psykiatrins
     33 psykiatrisk
     37 psykiatriska
      3 psykiatriskt
    116 psykisk
    174 psykiska
     61 psykiskt
      3 psykoaktiv
      8 psykoaktiva
      3 psykoaktivt
      1 psykoakustik
     16 psykoanalys
     28 psykoanalysen
      1 psykoanalysenexistentialismen
      8 psykoanalysens
      4 psykoanalytiker
      4 psykoanalytikern
     13 psykoanalytisk
     14 psykoanalytiska
      1 psykoanalytiskt
      2 psykodramaterapi
      1 psykodynamik
     15 psykodynamisk
      9 psykodynamiska
      1 psykodynamiskt
      1 psykoemotionella
     15 psykofarmaka
      1 psykofilosofi
      1 psykofysiologiska
     14 psykogen
      1 psykogena
      1 psykogent
      1 psykokirugi
      6 psykokirurgi
      3 psykokirurgiska
     13 psykolog
     12 psykologen
      1 psykologens
     19 psykologer
      1 psykologerkuratorer
      1 psykologerna
      1 psykologförbund
      1 psykologförbundet
      1 psykologhjälp
     25 psykologi
     17 psykologin
      5 psykologins
     33 psykologisk
     61 psykologiska
     10 psykologiskt
      1 psykologitermer
      1 psykologutbildningen
      2 psykometriskt
     13 psykomotorisk
      1 psykomotoriskt
      1 psykonauterna
      3 psykoneuroendokrinologi
      2 psykoneuroendokrinologin
      3 psykoneuroimmunologi
      2 psykoneuroser
      7 psykopat
     25 psykopaten
      5 psykopatens
     33 psykopater
      1 psykopaterna
     46 psykopati
      1 psykopatidrabbade
      1 psykopatikriterier
     14 psykopatin
      1 psykopatins
      4 psykopatisk
      6 psykopatiska
      1 psykopatitillståndet
      1 psykopatklasser
      4 psykopatologi
      6 psykopatologiska
      2 psykopats
    125 psykos
     39 psykosen
      4 psykosens
      1 psykosepisoder
    105 psykoser
      9 psykoserna
      2 psykosernas
      1 psykosers
      1 psykosexuella
      1 psykosexuellt
      1 psykosinsjuknandet
      1 psykoslindring
      1 psykoslindringen
      8 psykosocial
     20 psykosociala
      4 psykosocialt
      7 psykosomatisk
      7 psykosomatiska
      1 psykosomatiskt
      1 psykossjuka
      2 psykossjukdom
     11 psykossjukdomar
      1 psykossymptom
      2 psykossymtom
      1 psykostillståndet
      1 psykoterapeut
      2 psykoterapeuten
      4 psykoterapeuter
      3 psykoterapeutisk
      1 psykoterapeutiska
     40 psykoterapi
      1 psykoterapiernai
      1 psykoterapiform
      3 psykoterapiformer
      1 psykoterapikliniker
      1 psykoterapimetod
      5 psykoterapin
      1 psykoterapiorganisationen
     10 psykotisk
     33 psykotiska
      2 psykotiske
      1 psykotiskt
      8 psykotropkonvention
      4 pt
      2 pta
      2 ptah
      1 pterin
      2 pteronyssinus
      2 pth
      1 pthirus
      1 pthreceptordefekt
      3 ptk
      1 ptkäven
      1 ptkgenen
      1 ptoområdet
      1 ptos
      3 ptsd
      1 ptsta
     10 pu
      1 pubar
      1 pubchem
      1 pubertas
     12 pubertet
     62 puberteten
      1 pubertetsbedömning
      1 pubertetsbedömningen
      1 pubertetsrelaterade
      2 pubertetsutveckling
      3 pubertetsutvecklingen
      1 pubes
      3 pubescens
      2 pubesområdet
      1 pubesregionen
      2 pubiotomi
      4 pubis
      6 public
      2 publicera
      9 publicerad
      1 publiceradbr
     32 publicerade
     30 publicerades
      5 publicerar
      3 publiceras
     13 publicerat
      5 publicerats
      4 publicering
      2 publiceringen
      2 publiceringsbias
      1 publicitet
      1 publikation
      1 publikationen
      3 publikationer
      1 publiken
      1 publishers
      3 pubmed
      1 puckel
      2 puckelrygg
      1 pucoga
     13 puder
      1 puerperalpsykos
      1 puerperiets
      1 puerperium
      1 puerto
      1 puffa
      1 pukarispukeris
      1 pulex
      1 pulmicort
      3 pulmonalis
      1 pulmonalisangiografi
      2 pulmonalisklaffen
      1 pulmonalvenerna
      2 pulmonary
      3 pulmonell
      1 pulmonella
     33 puls
      3 pulsad
      1 pulsåderbråck
      1 pulsatilla
     11 pulsen
      2 pulsera
      3 pulserande
      1 pulserar
      1 pulsfrekvensen
      2 pulsmätning
      1 pulsoximetri
      2 pulsslag
      1 pulsus
     16 pulver
      3 pulverform
      1 pulverformiga
      1 pulverformigt
      4 pulverinhalator
      1 pulverinhalatorer
      1 pulverisera
      1 pulvermaterial
      1 pulvermetoden
      1 pulversoppor
      1 pulvinar
      2 pulvis
      4 pulvret
      1 pulvriserad
      1 pulvriserade
      1 pulvriserar
      3 pump
     13 pumpa
     11 pumpar
     20 pumpas
      1 pumpbehandling
      2 pumpen
      2 pumpförmåga
      1 pumpförmågan
      3 pumpfunktion
      1 pumpning
      1 punctura
      1 pund
      1 punding
      3 pung
      1 pungbråck
     21 pungen
      1 pungräv
      1 pungvred
      1 punkare
      1 punken
     13 punkt
     12 punkten
      1 punktens
     14 punkter
      1 punktera
      1 punkterad
      1 punkterar
      1 punktering
      5 punkterna
      2 punkternas
      1 punkterse
      3 punktion
      2 punktkombinationer
      1 punktmutation
      1 punktögon
      3 punktprevalens
      1 punktprevalensen
     11 punktskrift
      1 punktskriften
      3 punktskriftsbiblioteket
      1 punktskriftsbok
      1 punktskriftsböker
      1 punktskriftsmaskin
      2 punktskriftsskärm
      4 pupill
      1 pupilldilaterande
      8 pupillen
      1 pupillens
      5 pupiller
      1 pupillernas
      1 pupillförträngning
      2 pupillreaktion
      1 pupillreaktionerna
      2 pupillreaktionljusreflex
      1 pupillreflexen
      1 pupillsammandragningen
      1 pupillstorlek
      1 pupillutvidgning
      2 pupillvidgande
      3 puppa
      1 puppan
      1 puppor
      5 puppp
      2 puppstadiet
      1 puppstadium
      1 pure
      1 purgantia
      1 purgativ
      1 purified
      1 purin
      1 purinalkaloid
      1 purinderivat
      2 puriner
      1 purkinjefiber
      2 purkinjefibrer
      1 purkinjetrådar
      1 purkyn
      1 purpur
      5 purpura
      1 purpurae
      6 purpurea
      1 purpureafruitsjpgfrukter
      1 purpurfärgad
      2 purpurfärgade
      1 purpurröd
      1 purpurskatta
      1 purpursnäcka
      1 pus
      1 push
      3 pushup
      1 pushupbehå
      1 pushupbehåar
      1 pushupbh
      1 pushuptrend
      1 pusillus
      1 pussande
      3 pussel
      1 pusselbit
      1 pustertal
      1 putamen
      1 putamens
      1 putra
      2 putsa
      1 putta
      4 puumalavirus
      1 puumalaviruset
      1 puumalavirusets
      1 puuseppfrån
      1 puva
      1 pv
      5 pvåg
      4 pvågen
      1 pvågens
      1 pvågor
      1 pvärden
      1 pvcmattor
      1 pvk
      1 pvt
      1 pwcs
      1 pwr
      1 px
     11 pyelonefrit
      1 pyelonefriter
      1 pyelostomikateter
      1 pyemin
      1 pygméer
      2 pylonefrit
      4 pylori
      4 pylorus
      1 pylorusbihang
      1 pyloruskörtlar
      1 pylorusregionen
      3 pylorussfinktern
      1 pylos
      2 pyodermi
      1 pyogenes
      1 pyoryugi
      1 pyr
      1 pyraclostrobinazoxystrobin
      1 pyramidalcellers
      1 pyramidalcellsdendriterna
      1 pyramidbanan
      2 pyramiden
      1 pyramidloben
      1 pyran
      1 pyranring
      1 pyranringen
      2 pyrazinamid
      2 pyrenéerna
      1 pyretroidinsekticider
      1 pyrexi
      2 pyrodruvsyra
      3 pyrofosfat
      1 pyrofosfatkristaller
      1 pyrofosfatsynovit
      1 pyrogener
      1 pyrolys
      2 pyrolyseras
      1 pyromaner
      9 pyromani
      1 pyroteknik
      2 pyroxen
      4 pyroxener
      1 pyrroler
      2 pyrrolringar
      6 pyruvat
      1 pyrvin
      1 pytagoras
      1 pytagoréerna
      1 pythagoras
      1 pyttesmå
      1 pyuri
      1 pzl
      9 q
      1 q�
      2 qaly
      1 qalyan
      1 qassam
      1 qdeletion
      2 qdeletionsyndromet
     10 qfeber
     11 qi
      2 qigong
      2 qing
      2 qingdynastin
      1 qingzangjärnvägen
      1 qmärkt
      1 qmed
      1 qpotenser
      1 qrs
      2 qrskomplex
      6 qrskomplexet
      2 qt
      2 qtc
      2 qtsyndrom
      2 qttid
      2 qttiden
      1 quacken
      1 quacksalber
      2 quadrifolia
      1 quality
      1 quarantaine
      1 quarantena
      1 quattor
      1 quecksalber
      2 queen
      3 queensland
      1 quentinfängelset
      1 quervains
      1 query
      1 quesadillas
      2 questionnaire
      1 quetiapin
      1 quicks
      1 quincke
      1 quinckeödem
      2 quinoa
      1 quinquenervus
      2 quotient
      2 qvågen
      1 qvågsinfarkt
      1 qvarnström
      1 qvinligt
      1 qviström
     20 r
      1 ra
     11 rå
      9 råa
      2 raas
      1 raassystemet
      1 råbandsknopar
      1 rabarber
      1 rabarberliknande
      1 rabatter
      1 rabatteternell
      1 rabattväxt
      1 rabbla
      1 rabdomyo
      5 rabdomyolys
     29 rabies
      1 rabiesfall
      1 rabiesfria
      1 rabiesfritt
      1 rabiesimmunoglobuliner
      1 rabiesinfektion
      1 rabiessmitta
      1 rabiesvaccin
      1 rabiesvirus
      2 rabiesviruset
      3 racemat
      1 racemiskt
      1 racemosa
      1 rachmaninovs
     14 räcka
      1 räckbäcken
     49 räcker
      1 räckte
      1 raclopride
     82 rad
     41 råd
      1 rada
      1 råda
      9 rådande
      1 radarstationer
      1 rådata
     14 rädd
      1 rådda
     20 rädda
      1 räddade
      3 räddar
      1 räddare
      2 räddas
      5 räddat
      1 räddats
      3 rådde
      1 räddning
      1 räddningsarbetare
      1 räddningsarbetet
      1 räddningsinsatserna
      1 räddningsledare
      1 räddningsledaren
      3 räddningstjänst
      1 räddningstjänstbefäl
      1 räddningstjänsten
      1 räddningstjänstens
      1 räddningsverket
      2 raden
      1 råden
      3 rader
     42 råder
      8 rådet
      4 rådets
      1 rådfråga
      1 rådfrågas
      1 rådgivande
      1 rådgivare
      8 rådgivning
      1 radiala
      1 radiära
      1 radiärsymmetriska
      4 radiata
      5 radiation
      1 radicans
      3 radie
      1 radiella
      1 radien
      4 radikal
      1 radikala
      8 radikaler
      1 radikalerna
      1 radikalers
      1 radikalitet
      1 radikaloperation
      7 radikalt
      9 radio
      1 radioaktiv
     17 radioaktiva
      1 radioaktivitet
      1 radioaktiviteten
     14 radioaktivt
      2 radioapparater
      1 radiobiologi
      1 radiofarmaka
      1 radiofosfor
      1 radiofrekvensbehandling
      1 radiofrekvent
      2 radiofrequency
      5 radiofysik
      3 radiofysiken
      1 radiofysiska
      1 radiografi
      1 radiohead
      1 radiohitlåtar
      1 radioisotoper
      2 radiojod
      1 radiokirurgi
      1 radioligander
      1 radiolog
      1 radiologen
      1 radiologer
     15 radiologi
      1 radiological
      1 radiologin
      2 radiologisk
      5 radiologiska
      1 radiomottagning
      4 radionuklider
      1 radiophysique
      1 radiorör
      1 radiostörningar
      3 radioterapi
      2 radiotermoelektriska
      1 radiotrafiken
      1 radioutrustning
      1 radiovågor
      1 rädisor
      1 radium
      1 radiumhemmet
      2 radix
      7 rådjur
      1 rådjuren
      1 rådjurets
      7 radon
      1 radondöttrarnas
      1 radonets
      1 radongas
      1 radongashalten
      2 radonhalten
      1 radonkarbonatsmineralkällor
      1 radonrelaterade
      1 radonrisken
      2 råds
      1 räds
     82 rädsla
     20 rädslan
      7 rädslor
      1 rädsloreaktion
      1 rädsloreaktioner
      1 rädslorespons
      1 rädslorna
      1 raelians
      2 raffinerade
      1 raffinerat
      1 raffinering
      4 räfflad
      1 räfflade
      1 rafflesia
      6 råg
      1 ragad
      1 rågbröd
      1 raggarsträng
      1 raglande
      1 ragnar
      1 ragu
      1 ragú
      1 råguttaperka
      1 råguttaperkan
      1 raid
      1 raiders
      2 rail
      1 rain
      1 rajasthan
      3 rajayoga
      7 rak
     12 raka
      9 råka
      1 räka
      2 rakade
      3 råkade
      1 rakapparat
      1 rakapparaten
      1 rakar
      4 råkar
      1 rakare
      2 rakat
      5 råkat
      2 rakats
      5 rakborstar
      1 rakborstarna
      4 rakborste
      2 rakborsten
      1 rakborsthåret
      1 raketartilleriet
      1 raketdrift
      1 raketdysa
      1 raketer
      1 raketmotorer
      3 rakgel
      2 rakhyvel
      1 rakic
      6 rakit
      1 rakitis
      5 rakkniv
      2 rakknivar
      2 rakkniven
      1 rakknivsmärken
      3 rakkräm
      1 rakkrämer
      4 raklödder
     17 räkna
      2 räknade
      7 räknades
     39 räknar
      1 räknarens
      1 räknarna
    154 räknas
      7 räknat
      1 räknesten
      1 räknesvårigheter
     14 rakning
      5 räkning
      1 rakningen
      3 råkost
      1 råkostarianer
      2 råkostdieter
      1 rakprodukter
      1 raksasa
      2 rakskum
      1 raksträcka
     20 rakt
      1 rakta
      5 raktvål
      1 raktvålar
      3 rakvatten
      1 rålambsvägen
      1 raleigh
      1 rälerna
      1 ralf
      1 raloxifen
      2 ralph
      1 räls
      2 rälsen
      6 ram
      1 ramadan
      1 ramanujan
      1 ramarna
      1 ramas
      1 råmaterial
      1 ramdirektivet
      1 ramel
      8 ramen
      1 ramesseum
      1 råmjölk
      1 ramla
      1 ramlade
      2 ramlagar
      2 ramlar
      1 ramón
      2 rampfeber
      1 ramses
      1 ramsgate
      3 ramsor
      1 ramsystem
      1 ramverket
      2 rån
      1 rånat
      1 randar
      2 ränder
      1 randi
      2 randig
      2 randis
      3 randomiserad
      1 randomiserade
      1 randomiserades
      1 rånet
      1 rånförsök
      3 rang
      2 range
      1 ranglåg
      1 rangordnade
      1 rangordnas
      1 rankar
      1 rankat
      1 rann
      2 ränna
      1 rännan
      1 rännor
      1 ranstadsverket
      2 ränta
      1 räntebärande
      1 räntor
      1 ranunculus
     13 ranunkelväxter
      1 ranunkelväxternas
      1 ranviers
      1 råolja
      1 råoljebaserade
      2 rapa
      3 rapid
      1 rapning
      1 rapoport
      1 rappakalja
     29 rapport
     29 rapporten
     20 rapporter
     11 rapportera
      1 rapporterad
     32 rapporterade
     19 rapporterades
     10 rapporterar
      8 rapporteras
      4 rapporterat
     33 rapporterats
      7 rapportering
      4 rapporterna
      1 raps
      1 rapsbaggen
      1 rapsolja
      9 ras
      2 rasa
      2 rasade
      2 rasande
      1 rasanlag
      1 rasayana
      1 rasbiologi
      1 rasbiologiska
      4 rasen
      2 raser
      1 raseras
      4 raseri
      1 raserianfall
      1 raseriutbrott
      2 raserna
      1 rashad
      5 rashygien
      1 rashygienen
      2 rashygienens
      2 rashygieniska
      1 rashygieniskt
      1 rasilez
      1 rasism
      1 rasister
      1 raskatter
      2 raskt
      1 rasmussens
      2 rasoal
      1 rasoh
      6 rassel
      2 rassenhygiene
      2 rast
      1 rastar
      1 rasteori
      2 raster
      1 rastlöse
      3 rastlöshet
      1 rastlösheten
      1 rastlösthet
      2 rasttest
      2 rät
      3 räta
      1 ratade
      1 rätar
      2 rate
      1 rates
      1 ratificera
      1 ratificerade
      1 ratificerat
      2 rating
      1 ratio
      2 rational
      1 rationalisering
      1 rationalism
      3 rationell
      2 rationella
      2 rationellt
      1 ratt
      7 rått
    154 rätt
      8 råtta
     19 rätta
      5 råttan
      1 rättar
      1 rättare
      1 rättas
      1 råttblod
      1 rättegång
      1 ratten
     23 rätten
      1 rättesnöre
      1 rättfärdigar
      3 råttgift
      1 råtthonor
      3 rättighet
      1 rättigheten
     19 rättigheter
      1 rättigheterna
      1 rättning
     33 råttor
      2 råttorna
      2 råttors
      1 rättsfall
      1 rättsgenetik
      1 rättshandling
      3 rättshandlingar
      2 rättshandlingen
      1 rättsintyg
      1 rättsintyget
      1 rättskemi
      1 rättskrivning
      4 rättsläkare
      3 rättsläkaren
      2 rättslig
      1 rättsliga
      1 rättsligt
      9 rättsmedicin
      2 rättsmedicinalverket
      2 rättsmedicinalverkets
      1 rättsmedicinare
      4 rättsmedicinsk
      3 rättsmedicinska
      3 rättsodontolog
      1 rättsodontologen
      1 rättsodontologer
      1 rättsodontologi
      1 rättsodontologisk
      1 rättspraxis
      1 rättsprocesserna
      1 rättspsykiatisk
      4 rättspsykiatri
      6 rättspsykiatrin
      1 rättspsykiatrisk
      4 rättspsykiatriska
      1 rättsskandalen
      1 rättsstater
      2 rättssystem
      1 rättssystemet
      1 rättstraditionen
      1 rättsvårdande
      2 rättsväsendet
      2 rattus
      1 rättvisan
      1 rättvisande
      1 rättvisare
      1 raulin
      1 rav
      4 räv
      2 rävar
     11 råvara
      4 råvaran
      1 rävarnas
      9 råvaror
      2 råvarorna
      1 råvarornas
      1 råvarubörser
      1 råvarumarknaden
      2 rave
      1 ravens
      1 rävfett
      1 ravitch
      1 ravitchmetoden
      1 rävkaketräd
      1 rävskabb
      1 rävstatyett
      1 rävtörel
      3 raw
      1 rawfood
      1 ray
      1 rayban
      2 rayford
      1 raymi
      2 raymond
      2 rayner
      2 rayon
      1 raytheon
      6 rb
      1 rbcg
      1 rbgenen
      1 rctstudie
      1 rd
      2 rdi
      1 rditabell
      1 reabsoptionen
      1 reabsorberas
      7 reach
      2 reachsystemet
      5 reaction
      1 reactions
      1 reactor
      1 reading
      1 ready
      1 reagens
     42 reagera
      4 reagerade
      3 reagerande
     78 reagerar
      1 reageras
      1 reagerat
      3 reaginer
      1 reagintest
    106 reaktion
     31 reaktionen
      1 reaktionens
    124 reaktioner
      9 reaktionerna
      1 reaktionsförmåga
      1 reaktionskärlet
      1 reaktionskraft
      2 reaktionsmönster
      1 reaktionsprodukt
      1 reaktionstid
      1 reaktionsvägen
     11 reaktiv
     11 reaktiva
      1 reaktiverad
      1 reaktiveras
      2 reaktivering
      2 reaktivitet
      1 reaktiviteten
      1 reaktivt
      1 reaktor
      1 reaktorbränsle
      2 reaktorer
      3 real
      1 realgar
      1 realisera
      1 realiserad
      1 realisering
      2 realism
      2 realistisk
      3 realistiska
      2 realistiskt
      1 realitet
      1 realitetsprincipen
      2 reality
      1 realitysystem
      3 realtid
      1 realtidsavlyssning
      1 realtidsbevakningsteknologi
      1 realtidskonsultation
      1 realtidsvisning
      2 realtillgång
      1 realtillgångar
      1 realtime
      1 realvärdet
      2 reappraisal
      2 reassortment
      1 rebecka
      1 rebellen
      1 rebeller
      1 rebellsidan
      1 rebelsymbol
     19 recept
      3 receptarier
      3 receptbelagd
      6 receptbelagda
      8 receptbelagt
      1 recepten
      5 receptet
      1 receptets
      1 receptexpediering
      2 receptfri
     15 receptfria
      3 receptfritt
     12 receptor
     33 receptorer
      9 receptorerna
      1 receptorfamiljen
      1 receptormedierad
      1 receptormedierade
     10 receptorn
      1 receptorns
      1 receptors
      1 recessen
      2 recessiv
      4 recessivt
      5 recidiv
      4 recidiverande
      4 recip
      1 recipienten
      1 recitatör
      1 reckeweg
      1 reckitt
      2 recklinghausens
      1 reconstruction
      1 recorder
      1 records
      3 recruitment
      1 rectum
      1 rectus
      1 recycle
      3 red
     17 reda
      1 redaktionen
      1 redaktör
      1 redaktörsamma
    219 redan
      1 redden
      1 rede
      1 redi
      1 redigerad
      2 redigerats
      1 redlighet
      2 redlöst
      9 redo
      2 redogörelse
      5 redovisa
      2 redovisades
      1 redovisar
      1 redovisas
      2 redovisats
      1 redovisning
      1 redoxreaktion
      1 redressering
     17 redskap
      1 reduce
     31 reducera
      7 reducerad
      7 reducerade
      2 reducerades
      2 reducerande
     14 reducerar
     16 reduceras
      4 reducerat
      2 reducerats
      3 reducering
      1 reduceringen
      1 reductil
      2 reduction
      1 �reduktas
      5 reduktion
      1 reduktionen
      1 reduktionism
      1 reduktionsdelning
      2 reduktionsmissbildning
      1 reduktiv
      1 reed
      1 reelermössensknockoutmössens
      6 reelin
      1 reella
      1 reellt
      1 reevaluation
      1 ref
      1 refereegranskning
      3 references
      1 referenceshttpkisekijsppolopolyjsplsvda
      6 referens
      2 referensdata
      1 referenselektrod
     22 referenser
      1 referenserna
      1 referensgruppen
      1 referensintervall
      1 referenslista
      1 referensområde
      1 referenspunkt
      1 referenspunkter
      1 referensram
      1 referenssignal
      2 referensvärde
      1 referensvärden
      3 referensvärdena
      1 referensvärdenaför
      3 referera
      1 refererad
      2 refererade
     17 refererar
      4 refereras
      1 refererats
      1 reflektera
      2 reflekterade
      5 reflekterande
      5 reflekterar
      5 reflekteras
      2 reflekterat
      2 reflektion
      1 reflektioner
     13 reflex
     14 reflexen
      2 reflexens
      7 reflexer
      3 reflexerna
      2 reflexionsgoniometern
      1 reflexiva
      1 reflexmässig
      1 reflexmässiga
      1 reflexmässigt
      1 reflexmönster
      1 reflexologi
      1 reflexsammandragning
      1 reflexstyrd
      1 reflexutvecklingen
      1 reflexzonterapi
      5 reflux
      3 refluxesofagit
      1 reform
      1 reformen
      2 reformer
      1 reformliv
      1 refusal
    172 regel
      1 regelbrott
     15 regelbunden
      1 regelbundenhet
     44 regelbundet
     21 regelbundna
      1 regelmässig
      1 regelmässiga
      5 regelmässigt
      4 regeln
      1 regelrätta
      1 regelsystemen
      1 regelsystemet
      3 regelverk
      2 regelverket
      1 regementen
      1 regeneration
      1 regenerera
      1 regenererande
      1 regenereras
      1 regenerering
      7 regering
      5 regeringar
     21 regeringen
      1 regeringens
      1 regeringriksdag
      1 regerings
      1 regeringschefer
      1 regeringscheferna
      1 regeringsnivå
      1 regeringspolicyer
      1 regeringsproposition
      1 regeringsrätten
      1 regeringsuppdrag
      1 reggaeton
      5 regi
      1 regimen
      3 region
      5 regional
      8 regionala
      1 regionalkontor
      1 regionalt
      8 regionen
      2 regionens
     27 regioner
      3 regionerna
      1 regionkliniken
      1 regionkliniker
      1 regionsjukhus
      1 regionsjukhusen
      1 regionsjukhuset
      1 regionsklinik
      1 regisserad
      5 register
      2 registerbrott
      1 registerstudier
      1 registration
     12 registrera
      9 registrerade
      2 registrerades
     13 registrerar
     24 registreras
      4 registrerat
      1 registrerats
      8 registrering
      3 registreringen
      1 registreringsförmåga
      1 registreringsmetoder
      1 registreringsnatten
      1 registreringsprocedurer
      2 registreringstiden
      1 registreringstvånget
      1 registreringsutrustning
      1 registreringsutrustningen
      2 registret
      3 reglemente
      4 reglementen
     38 regler
     31 reglera
     11 reglerad
      3 reglerade
      2 reglerades
      6 reglerande
     35 reglerar
     28 regleras
      6 reglerat
      2 reglerats
      1 reglerbar
     22 reglering
      2 regleringar
     13 regleringen
      1 regleringskraften
     13 reglerna
      8 regn
      1 regna
      1 regnar
      1 regnbåge
      2 regnbågshinna
      2 regnbågshinnan
      1 regnbågshinnaniris
      2 regnbågshinneinflammation
      1 regnform
      1 regniga
      1 regnperioden
      2 regnskogen
      1 regntiderna
      1 regnvatten
      1 regress
      3 regression
      1 regular
      1 regulatorisk
      1 regulatorn
      1 regulatory
      1 reguljärt
      2 rehab
      1 rehabhund
      2 rehabilitera
      1 rehabiliterar
      1 rehabiliteras
     31 rehabilitering
      6 rehabiliteringen
      2 rehabiliteringsarbete
      1 rehabiliteringsåtgärd
      1 rehabiliteringsinsatser
      1 rehabiliteringsinsatserna
      1 rehabiliteringskostnader
      1 rehabiliteringsmedicin
      1 rehabiliteringsmetoder
      1 rehabiliteringsperioden
      1 rehabiliteringsprojekt
      1 rehabiliteringsträning
      1 rehållning
      1 rehydrex
      1 reich
      1 reichsführerss
      1 reiki
      1 reil
      1 reisseissenmuskler
      3 reiters
      1 rejäl
      3 rejäla
      1 rejält
      1 rejektion
      1 rejektvatten
      2 rejuvelac
      3 reklam
      1 reklamen
      1 reklamfilm
      1 reklamföra
      1 reklamkampanjer
      1 reklampionjären
      1 reklamstoppet
      3 rekombinant
      2 rekombinanta
      1 rekombination
      1 rekomenderas
     12 rekommendation
      4 rekommendationen
     13 rekommendationer
      5 rekommendationerna
      7 rekommendera
      5 rekommenderad
     12 rekommenderade
      4 rekommenderades
     40 rekommenderar
    113 rekommenderas
      9 rekommenderat
      1 rekommenderats
      1 rekompressionsbehandling
      2 rekonstruera
      2 rekonstruerade
      7 rekonstruktion
      1 rekonstruktioner
      1 rekonstruktionskirurgi
      6 rekonstruktiv
      1 rekonstruktiva
      1 rekord
      4 rekordbok
      1 rekordnotering
      2 rekreation
      1 rekreationella
      3 rekreationellt
      1 rekreationen
      1 rekreationsanläggningar
      2 rekreationsdrog
      1 rekreationsdykare
      1 rekreationskonsumenter
      2 rekreationskonsumtion
      2 rekryterar
      2 rekrytering
      5 rektal
      4 rektala
      3 rektalt
      1 rektangel
      1 rektangulär
      2 rektoskopi
      2 rektum
      1 rekvisita
      1 relä
      1 relästation
      2 related
      4 relatera
     12 relaterad
     20 relaterade
      1 relaterades
      2 relaterar
      4 relateras
     20 relaterat
      1 relaterats
     31 relation
      1 relationell
      1 relationella
      9 relationen
     37 relationer
      2 relationerna
      2 relationsproblem
      1 relationsskapande
      3 relativ
     13 relativa
      1 relativisera
      1 relativiserar
    180 relativt
      1 relau
      1 relaxation
      1 relaxering
      1 relaxin
      1 releaseinhibiting
      1 relegering
      1 releterade
      1 relevance
      2 relevans
      1 relevansen
     11 relevant
      9 relevanta
      1 reliabilitet
      1 reliabiliteten
      1 reliability
      1 relief
      8 religion
      2 religionen
     13 religioner
      4 religionerna
      1 religioners
      1 religionsgränserna
      1 religionsgrundaren
      1 religionshistoriker
      1 religionspolis
      1 religionsvetenskapligt
     11 religiös
     35 religiösa
      4 religiöst
      1 relikskrin
      1 relikt
      1 reliktro
      5 rem
      1 remdrivna
      1 remedia
      1 remember
      2 remifentanil
      1 remifentanilanestesi
      1 remineralisationshastighet
      1 reminyl
      1 reminylgalantamin
      2 remiss
      1 remissförfarande
      5 remission
      1 remittent
      3 remittera
      1 remitterar
      3 remitteras
      1 remitting
      1 remlika
      2 remmar
      1 remodellerade
      1 remover
      1 remperiod
      2 remsa
      3 remsan
     15 remsömn
      8 remsömnen
      1 remsömntiden
      1 remsor
      1 remsorna
     61 ren
     36 rena
      4 renade
      4 renal
      1 renalt
      6 renande
      4 renar
      1 renare
      2 renarna
     18 renas
      2 renässans
     10 renässansen
      1 renässansmänniskor
      1 renaste
      1 renat
      1 renderar
      1 rendezvouz
      1 rene
      4 rené
      5 renens
      1 renframställa
      1 rengjord
      2 rengjorda
      1 rengjorde
      2 rengjordes
      1 rengjort
      1 rengjorts
      4 rengör
     17 rengöra
      1 rengörande
      3 rengöras
     31 rengöring
      1 rengöringslösningar
     19 rengöringsmedel
      1 rengöringsproblem
      1 rengöringsprocessen
      1 rengöringsprodukter
      2 rengörs
      1 renhållning
      1 renhållningsarbete
      4 renhet
      1 renhjärta
      1 renhjordarna
      8 renin
      1 reninangiotensin
      1 reninangiotensinaldosteronsystemet
      5 reninangiotensinsystemet
      1 reninfrisättning
     15 rening
      6 reningen
      1 reningsgrad
      1 reningsprocess
      1 reningsprocessen
      1 reningssteget
      3 reningsverk
      1 reningsverken
      1 reningsverkens
      5 reningsverket
      2 reninhämmare
      1 reninhämning
      1 renis
      2 renläriga
      1 renlevnad
      1 renlevnads
      5 renlighet
      1 renodlad
      4 renodlade
      1 renodlades
      1 renografi
      1 renoveras
      1 renovering
      1 renparasiten
      4 renrum
      7 rensa
      1 rensad
      2 rensar
      2 rensas
      1 rensat
      1 renset
      1 rensgaller
      2 rensgallret
      1 renshaw
      1 renskinn
      1 renskötare
      2 renskötselområden
      1 renskötselområdena
      1 renslakt
      1 renströmska
      4 renstyng
      3 renstynget
      2 renstyngets
      1 renstyngsfluga
      1 renstyngsflugan
     88 rent
      3 rentav
      1 rentutav
      1 reoviridae
      4 rep
      1 repair
      3 reparation
      1 reparationsförmåga
      1 reparationskostnader
      1 reparationsmateriel
      1 reparationssystem
      5 reparera
      1 reparerar
      4 repareras
      1 repellera
      1 repens
      1 repeteras
      1 repetetiva
      1 repetitiv
      3 repetitiva
      5 repetitivt
      1 replik
      3 replikation
      1 replikationscykel
      1 repliker
      1 replikera
      2 replikerar
      1 replikeras
      1 replikerbar
      1 replikering
      2 repolarisation
      2 repolarisationen
      2 repolarisering
      5 repor
      1 reportern
      1 reportrar
      1 repositioning
      9 representanter
      4 representation
      1 representationen
     10 representationer
      2 representationerna
      2 representativ
      2 representativa
      1 representativt
      5 representera
      5 representerad
      6 representerade
      1 representerades
     16 representerar
      8 representeras
      1 representerat
      1 repression
      1 reprocessing
      3 reproducera
      1 reproducerade
      1 reproducerande
      2 reproducerar
      3 reproduceras
      1 reproducerbar
      1 reproducerbara
     10 reproduktion
      2 reproduktionen
      1 reproduktionsapparaten
      1 reproduktionsförmågan
      2 reproduktionsmedicin
      1 reproduktionsmekanismer
      4 reproduktionsorgan
      1 reproduktionssättet
      1 reproduktionssystem
      2 reproduktionssystemet
      5 reproduktiv
      5 reproduktiva
      1 repslagning
      3 reptåliga
     10 reptiler
      1 reptition
     10 republiken
      1 repulsion
      1 repulsiva
      1 requiem
     11 resa
      1 resacetofenon
      6 resan
      7 resande
      1 resår
      1 resårer
     14 research
      1 researchers
      1 resebagaget
      2 reseetui
      3 resektion
      1 resenärer
      9 reser
      1 reserpin
      1 reservaten
      1 reservdroger
      1 reserver
      1 reserverad
      2 reserverade
      1 reserverna
      2 reservkapacitet
      2 reservmediciner
     11 reservoar
      6 reservoaren
      1 reservoirer
      1 resetidningen
      1 resetransport
      1 resevaccinationer
      1 residual
      1 residualschizofreni
      1 resisens
      1 resistance
      7 resistans
      5 resistansen
      1 resistansmekanismer
      2 resistena
     83 resistens
      6 resistensen
      1 resistensfrekvensen
      4 resistensgener
      1 resistensgenerna
      2 resistensmekanism
      2 resistensproblem
      1 resistensproblemet
      4 resistensspridning
      2 resistensspridningen
      6 resistensutveckling
      1 resistensutvecklingbehandlingstiden
      1 resistensutvecklingen
     11 resistent
     40 resistenta
      1 resistentare
      2 resistin
      3 resistorer
      1 resmål
      1 resmålet
      1 resningen
      5 resolution
      1 resolutioner
      1 resonance
      4 resonans
      3 resonansen
      4 resonanser
      1 resonansformer
      2 resonansfrekvens
      1 resonansfrekvenser
      1 resonanskrets
      2 resonanslåda
      1 resonanslådan
      1 resonansmönster
      1 resonansrummet
      1 resonansstrukturer
      5 resonanstomografi
      2 resonemang
      1 resonemangen
      1 resonemanget
      4 resonera
      1 resonerar
      1 resonsstrukturer
      9 resor
      1 resorbera
      3 resorberas
     10 resorberbara
      1 resorberingen
      6 resorcinol
      1 resorna
      3 resource
      5 resp
      1 respekt
      1 respekterad
      1 respekteras
      1 respektfullt
    127 respektive
      1 respektlös
      1 respirabla
      5 respiration
      1 respirationsfysiologi
      1 respirationsfysiologin
      1 respirationshistologi
      1 respirationssystemet
      1 respirationsvägarna
     10 respirator
      1 respiratorbehandlas
      3 respiratorbehandling
      1 respiratorbehandlingcpap
      2 respiratorbehandlingen
      6 respiratorer
      1 respiratorerna
      1 respiratorii
     22 respiratorisk
      3 respiratoriska
      3 respiratoriskt
     10 respiratorn
      1 respiratorvård
      3 respiratory
      1 respironics
      1 respondenten
      1 respondenter
     22 respons
      6 responsen
      4 responser
      1 responsiva
      3 responsprevention
      1 responspreventionen
      1 responssyndrom
      1 responstid
      5 rest
      3 restaurang
      1 restaurangen
     11 restauranger
      1 restaurera
      1 restaurerades
      6 reste
     39 resten
      1 restenos
     17 rester
      9 resterande
      4 resterna
      1 restes
      1 restmetaboliter
      3 reston
      2 restprodukt
      6 restprodukter
      2 restprodukterna
      1 restriction
      8 restriktioner
      1 restriktionerna
      8 restriktiv
      4 restriktiva
      2 restriktivt
      1 restskada
      3 resttillstånd
      4 restylane
    168 resultat
     44 resultaten
     70 resultatet
      1 resultatets
      1 resultatlösa
     17 resultera
     16 resulterade
      2 resulterande
     44 resulterar
      5 resulterat
      2 resurs
      1 resursbegränsade
      1 resursbrist
      1 resurscentra
     18 resurser
      1 resursstarka
      1 resurssvaga
      1 resvanor
      3 retande
      6 retar
      8 retardation
      1 retardering
      1 retbara
      1 retbarheten
      2 retention
      2 rethosta
      1 retia
      2 reticularis
      1 reticulata
      1 reticulosa
      1 reticulum
      1 retiklet
     11 retikulära
      1 retikulocyter
      4 retina
      2 retinal
      1 retinasjukdom
      1 retinitis
     10 retinoblastom
      1 retinoblastomen
      2 retinoblastomprotein
      1 retinol
      1 retinopathy
      2 retirerar
      1 retledning
      1 retledningshinder
      1 retledningssystem
      1 retledningsystem
      1 retliga
      1 retlighet
      7 retning
      2 retningarna
      2 retningen
      1 retoriken
      2 retraining
      1 reträttmarsch
      1 retriever
      1 retrievrar
      2 retrograd
      1 retrokänsla
      3 retrospektiv
      3 retrospektiva
      2 retrovirus
      1 retroviruset
      4 retts
      2 returfiber
      2 returfiberbaserade
      1 returpapper
      2 returslam
      2 retzius
      1 reumatiker
      8 reumatisk
      8 reumatiska
     13 reumatism
     10 reumatoid
      1 reumatologen
      2 reumatologisk
      2 reumatologiska
      1 réunion
      1 reuse
      1 reuteri
      1 reuters
      9 revben
      7 revbenen
      1 revbenets
      1 revbensbåge
      1 revbensbågen
      1 revbensbrosken
      1 revbensbrott
      1 revenue
      1 reversal
      1 reverse
      1 reversera
      6 reversibel
      1 reversibilitetstest
      2 reversibla
      1 reviderades
      1 reviderat
      3 reviderats
      3 revidering
      7 review
      1 reviews
      1 revirstrider
      1 revised
      2 revisionen
      1 revisioner
      1 revolt
      1 revoltbenägen
      7 revolutionen
      2 revolutionerade
      1 revolutionerades
      1 revolutionerat
      2 revor
      1 revorm
      3 revsmörblomma
      1 revsmörblommans
      1 rexona
      4 reynolds
      1 rf
      1 rfablation
      1 rfc
      1 rfel
      1 rfhl
      1 rform
      2 rformen
      2 rfsl
      2 rfsu
      1 rgrm
     16 rh
      1 rhabdomyom
      2 rhabdomyosarkom
      2 rhabdoviridae
      1 rhabdovirus
      1 rhabidoviridae
      1 rhd
      1 rhenium
      1 rheo
      2 rhesus
      1 rhesusantigen
      1 rhesusapan
      1 rhesusapor
      2 rhesusfaktorn
      1 rhett
      1 rheuma
      1 rhinit
      1 rhinkompatibilitet
      1 rhino
      1 rhinotillexomani
     14 rhinovirus
      5 rhinoviruset
      1 rhinovirusförkylningar
      1 rhinovirusinfektionens
      1 rhizobium
      2 rhizomorfer
      1 rhizomorferna
      1 rhnegativ
      1 rhnegativt
      1 rhodesiense
      1 rhododendron
      1 rhododendronarter
      1 rhoos
      1 rhpositiv
      4 rhsystemet
      1 rhynchophthirina
      5 ribavirin
      1 ribbade
      1 ribes
      1 ribonukleas
      1 ribonukleinsyra
      1 ribonukleinsyran
      1 ribos
      4 ribosomen
      8 ribosomer
      2 ribosomerna
      1 ricardo
     17 richard
      1 richelieu
      1 richet
      3 ricinolja
      1 ricinus
      1 ricinus]
      1 rickettsia
      1 rickettsiabakterier
      1 rickettsibakterier
      1 rickettsier
      1 ricky
      1 rico
      1 rid
      1 ridande
      1 ridbågarna
      1 riddarmusseron
      1 riddarsporresläktet
      1 riddjur
      2 rider
      1 ridge
      1 ridhjälmen
      1 ridley
      2 ridväg
      1 riesengebirge
     12 rifampicin
      6 rifampin
      1 rifamycin
      1 rige
      1 rigga
      1 riggad
      1 right
      1 rights
      2 rigiditet
      1 rigidula
      1 rigidus
      1 rigmor
      3 rigoröst
      1 rigveda
     20 rik
     14 rika
      3 rikare
      2 rikaste
      3 rikedom
      7 riket
      4 rikets
      9 riklig
      4 rikliga
      1 rikligare
     11 rikligt
      1 riksangelägenhet
      1 riksansvar
      1 riksbanken
      1 riksbanker
      1 riksbekant
      3 riksdag
      2 riksdagen
      1 riksdagsledamöter
      6 riksförbund
      5 riksförbundet
      1 riksförbunds
      2 riksföreningen
      1 riksinstruktören
      1 rikslikare
      1 riksomfattande
      2 riksorganisation
      1 riksperoner
      1 rikspolisstyrelsen
      1 rikspolisstyrelsens
      1 riksreglemente
      1 rikssjukhus
      1 riksstaden
      1 rikssvenskt
      1 riksväg
      1 riksvapnet
      5 rikt
      7 rikta
     10 riktad
     13 riktade
      1 riktades
     18 riktar
     12 riktas
      8 riktat
      1 riktats
      9 riktig
     11 riktiga
     28 riktigt
      1 riktlinje
     24 riktlinjer
      6 riktlinjerna
     24 riktning
     11 riktningar
      3 riktningen
      1 riktvärde
      1 riktvärden
      1 riktvärdet
      1 rima
      2 rimantadin
      5 rimlig
      3 rimliga
      1 rimligen
      4 rimligt
      1 rimma
      1 rimmad
      1 rimmande
      3 rinca
      1 rinderpest
      1 rinexin
     15 ring
     11 ringa
      1 ringaktning
     10 ringar
      2 ringarna
      1 ringbärande
      2 ringborg
      1 ringborgs
      1 ringbrosk
      1 ringbrosket
      2 ringbroskkannbroskmuskeln
     11 ringen
      3 ringer
      1 ringeracetat
      2 ringfingret
      1 ringformad
      1 ringformat
      1 ringla
      2 ringlar
      1 ringmärkning
      1 ringmaskarna
      1 ringmuskel
      2 ringmuskeln
      2 ringmuskler
      1 ringningar
      1 ringorm
      1 ringstadium
      1 ringstruktur
      3 rinit
     10 rinna
     18 rinnande
     11 rinner
      1 rinniga
      1 rinnsnuva
      1 rinofaryngit
      1 rinokonjunktivit
      1 rinologi
      1 rinologin
      1 rinorré
      1 rinosinuit
     20 ris
      1 risdrycker
      1 risets
      1 risi
    278 risk
      1 riskabel
      6 riskabelt
      1 riskabla
      1 riskan
      1 riskanalys
      3 riskbedömning
      8 riskbedömningar
      1 riskbedömningen
      1 riskbefolkningen
      2 riskbeteende
      4 riskbruk
    325 risken
     51 risker
      9 riskera
     38 riskerar
     33 riskerna
     13 riskfaktor
     47 riskfaktorer
      4 riskfaktorerna
      4 riskfaktorn
      2 riskfri
      3 riskfritt
      1 riskfyllda
      2 riskfyllt
      2 riskgrupp
     12 riskgrupper
      1 riskgrupperna
      1 riskhomeostas
      1 riskhomeostasteorin
      1 riskkällor
      1 riskkvoterna
      1 risknivå
      1 risknivån
      4 riskökning
      1 riskökningen
      2 riskområden
      1 riskorgan
      2 riskorna
      2 riskpatienter
      1 riskpersoner
      1 risksänkare
      3 risktagande
      1 risktagandet
      1 risktillfället
      2 riskuppfattning
      1 riskuppskattning
      1 riskvärderingar
      1 riskzon
      8 riskzonen
      1 risodling
      1 risomeren
      1 rispades
      1 rispas
      3 risperidon
      3 risperidone
      1 rispningar
      2 rispor
      1 risrätter
      1 risus
      5 rita
      1 ritade
      1 ritalin
      7 ritas
      1 ritat
      2 riter
      3 ritual
      3 ritualen
     16 ritualer
      3 ritualerna
      2 ritualistisk
      4 rituell
      5 rituella
      1 rituellt
      3 rituximab
      1 riv
      2 riva
      1 rivas
      2 rivastigmin
      4 river
      1 rivieran
      3 rivning
      1 rivningen
      1 rivningsarbetare
      1 rivningsarbete
      1 rivningsarbeten
      1 rivningstillstånd
      1 rivsår
      5 rls
     14 rna
      1 �rna
      1 rnamolekylen
      3 rnapolymeras
      1 rnapolymeraset
      1 rnaritningar
      2 rnasyntesen
      1 rnatyp
      6 rnavirus
      4 rns
      1 ro
      1 roa
      1 roanläggning
      1 roar
      1 rob
     22 robert
      1 roberto
      1 roberts
      1 robertsonfenomen
      2 robin
      2 robles
      3 robomemo
      1 robot
      1 robotar
      1 robotassisterade
      3 robust
      1 rochas
      6 rock
      1 rockar
      1 rockarnas
      1 rockartister
      1 rocken
      1 rocketbelt
      1 rockgrupper
      1 rockikonen
      1 rockkonsert
      1 rockland
     36 röd
    118 röda
      4 rödaktig
      1 rödaktiga
      1 rödaktigarosa
      1 rödaktigt
      1 rödalg
      1 rödalgerna
      1 rödare
      1 rödblåfärgade
      4 rödbrun
      2 rödbruna
      1 rödbrunaktiga
      2 rödbrunt
      1 rödceder
      1 rodd
      2 rodenticid
      1 rodeos
      1 rödfärga
      1 rödfärgad
      1 rödfärgade
      1 rödfärgat
      1 rödfläckig
      1 rödflammig
      1 rödflammiga
      1 rödflammigt
      1 rödgul
      2 rödgula
      1 rödkål
      1 rödlila
      2 rödlista
      4 rödlistad
      1 rödmaneter
      1 rödmaneterna
      1 rodna
     32 rodnad
      1 rodnade
      1 rödnade
      6 rodnaden
      4 rodnader
      3 rodnande
      4 rodnar
      2 rodnat
      1 rodolfo
      1 rodopsin
      1 rödräv
      1 rödräven
      1 rodríguez
      1 rödrosa
      1 rödsjuka
      2 rödsot
      1 rödsprit
      2 rödviolett
      1 rödvioletta
      1 rödvit
      4 rofecoxib
      1 roger
      2 rogivande
      1 rohm
      1 roine
      1 röja
     14 rök
     30 röka
      5 rökande
      1 rökandet
     19 rökare
      1 rökaren
      1 rökares
      1 rökarna
      2 rökas
      6 rökavvänjning
      1 rökavvänjningsprogram
      2 rökbad
      2 rökbastu
      2 rökbastun
      1 rökdetektorer
      1 rökdoften
      7 rökdon
      1 rökdonen
      1 rökdonet
      2 rökelse
      1 rökelsebehållaren
      1 rökelsebrännaren
      1 rökelsefatet
      1 rökelseritualer
      1 rökelsestickor
      6 röken
     14 röker
      8 rökförbud
      2 rökförbudet
      1 rökfrekvensen
      2 rökgång
      1 rökgaserna
      1 rökgasrening
      2 rökiga
      2 rokitansky
      2 rökmaterialet
    111 rökning
      1 rökningar
      7 rökningen
      2 rökningens
      1 rökningsmotståndares
      3 rökrör
      4 röks
      1 röksignaler
      1 rökskador
      3 rökstopp
      5 rökt
      2 rökta
     11 rökte
      5 röktes
      2 rökts
      1 röktsaltat
      1 rökvanor
      4 rolf
      5 rolfing
    107 roll
      3 rollator
      5 rollatorer
      5 rollatorn
      1 rollatortätaste
      1 rollekar
      4 rollen
      2 roller
      1 rollerna
      2 rollfigur
      2 rollon
      1 rolls
      5 rollspel
      1 rollvibration
     22 rom
      9 roman
      2 romanen
      2 romaner
      1 romanserien
      2 romanska
      1 romansvit
      1 romantik
      2 romantiken
      1 romantiserad
      1 romantiserades
      1 romantiserar
      3 romantiska
      1 romare
      1 romaren
      6 romarna
      3 romarnas
      1 romarrike
      3 romarriket
      1 romartid
      1 romartiden
      2 rombiska
      1 romeo
      2 romer
      1 romero
      6 romersk
     10 romerska
      2 romerske
      2 romerskkatolska
      1 rommel
      1 roms
      3 ron
      7 rön
      2 ronald
      1 rondeller
      1 rondo
      1 rondskål
      1 rönen
      3 ronki
      1 ronnie
      1 ronsard
      1 rönt
      1 röntga
     19 röntgen
      1 röntgenanalys
      2 röntgenapparaten
      1 röntgenapparatur
      1 röntgenavdelningar
      5 röntgenbild
      1 röntgenbilden
      9 röntgenbilder
      1 röntgenbilderna
      2 röntgenbildtagning
      1 röntgenfilmer
      1 röntgenfotografier
      1 röntgenfynd
      2 röntgengenomlysning
      1 röntgeninformationssystem
      1 röntgeninstitut
      1 röntgenkliniken
      5 röntgenkontrastmedel
      4 röntgenkristallografi
      1 röntgenkristallografin
      2 röntgenkristallografisk
      2 röntgenläkaren
      1 röntgenlaser
      1 röntgenmöte
      1 röntgenografik
      1 röntgenologisk
      2 röntgenologiska
      4 röntgenrör
      1 röntgenrum
      2 röntgensjuksköterskor
      1 röntgenspektrografi
      1 röntgenspektroskopi
      2 röntgenstrålar
      1 röntgenstrålarna
      1 röntgenstrålarnas
      2 röntgenstråldos
     19 röntgenstrålning
      2 röntgenstrålningen
      4 röntgenstrålningens
      1 röntgenstrålningsområdet
      1 röntgenundersöka
     22 röntgenundersökning
      7 röntgenundersökningar
      1 röntgenundersökningen
      1 röntgenvåglängder
      1 roosevelt
      6 rop
      1 ropade
      1 ropar
      1 ropet
    123 rör
     51 röra
     19 rörande
      1 röras
      4 rörben
      1 rörbenen
      1 rörbenens
      1 rörblad
      1 rörbladens
      6 rörde
     44 rörelse
      3 rörelseanalys
      1 rörelseanalyser
      1 rörelseanalyssystem
      3 rörelseapparat
      4 rörelseapparaten
      1 rörelsecentrum
      4 rörelseenergi
      1 rörelseenergin
      1 rörelsefunktion
      1 rörelsefunktionen
      1 rörelsehandikapp
      2 rörelsehinder
      1 rörelsehindrade
      1 rörelseinskränkningar
      2 rörelsekonst
      1 rörelsekonstnärer
      1 rörelsekraft
      1 rörelsekraften
      1 rörelsemoment
      6 rörelsemönster
      1 rörelsemönstret
     22 rörelsen
      1 rörelsenerv
      1 rörelsens
      1 rörelseövningar
      1 rörelseprogram
     74 rörelser
      1 rörelserädsla
      1 rörelseriktningar
      9 rörelserna
      5 rörelserubbningar
      1 rörelserutinen
     10 rörelsesjuka
      1 rörelsesjukdom
      1 rörelsesjukdomar
      1 rörelsestörning
      1 rörelsestörningar
      1 rörelsestörningarna
      4 rören
      1 rörens
      3 röret
      1 rörformade
      3 rörformat
      1 rörformiga
      2 rörformigt
      1 rörinstallationer
      2 rörledningar
     10 rörlig
     17 rörliga
      1 rörligare
     16 rörlighet
      4 rörligheten
      2 rörligt
      1 rörlika
      2 rörs
      1 rörsegement
      1 rörsegmenten
      1 rörsegmentens
      4 rört
      1 ros
      1 rós
     23 rosa
      1 rosace�
      2 rosafärgade
      1 rosalie
      1 rosatonad
      1 rosdahl
      1 rose
      1 rosemary
      2 rosen
      1 rosenblad
      1 rosenborgs
      1 rosenflockelssläktet
      1 rosenhall
      1 rosenhans
      1 rosenkvitten
      1 rosenlager
      1 rosenlundsbadet
      4 rosenmetoden
      1 rosenmetodens
      1 rosenolja
      1 rosenrörelsepedagoger
      1 rosensköna
      1 rosenterapeuten
      3 rosenterapeuter
      1 rosenthal
      1 roses
      1 rosett
      1 rosettformigt
      2 roseus
      7 rosfeber
      1 roslagen
      1 roslagssjukan
      1 rosling
      1 rosmarin
      1 rosmarinus
      1 rosor
      1 rossellini
      1 rössner
     24 röst
      1 rösta
      2 röstade
      1 röstades
      1 röstalstring
      1 röstansträngning
      1 röstanvändning
      2 röstanvändningen
      1 röstbehandling
      1 röstbeteende
      3 röstbeteendet
     47 rösten
      2 röstens
     19 röster
      4 rösterna
      1 rostfärgat
      2 rostfria
      8 rostfritt
      1 röstfunktion
      1 röstgenerator
      1 rösthallucination
      3 rösthallucinationer
      1 rostiga
      1 röstigenkänning
      1 röstkälla
      5 röstkällan
      2 röstkvalitet
      2 röstkvaliteten
      2 röstläge
      1 röstlägen
      1 rostning
      1 röstningsförfarandet
      1 röstpåverkan
      7 röstproblem
      4 rösträtt
      2 röstregistret
      4 röstrubbning
      3 röstrubbningar
      1 rostskyddsfärg
      1 rostskyddspigment
      1 röstspringa
      8 röstspringan
      1 röststörning
      7 röststörningar
      1 röststörningarna
      7 röststyrka
      7 röststyrkan
      1 rostsvampar
      1 röstsyntes
      1 röstsyntetiserare
      3 röstteknik
      1 rösttekniken
      1 rösttekniktips
      6 röstterapi
      4 rösttrötthet
      2 röstventil
      1 röstyrken
      1 rosväxter
      1 rosväxterna
      9 rot
      2 rota
      1 röta
      2 rotad
      1 rötades
      1 rotanlaget
      3 rotation
      2 rotationen
      1 rotationer
      1 rotationsriktning
      1 rotatorier
     15 rotavirus
      2 rotavirusinfektion
      1 rotavirusinfektioner
      1 rotaviruspartikel
      1 rotavirusvaccin
      1 rotavirusvaccination
      2 rotbehandling
     14 roten
      1 rotens
      2 rotera
      1 roterad
      1 roterade
      1 roterades
      2 roterande
      5 roterar
      3 rotfrukter
      1 rotfyllda
      1 rotfyllning
      1 rotfyllningen
      1 rotfyllningsmetoden
      1 rötgas
      4 rötgasen
      1 rötkammare
      1 rotkanaler
      1 rotkanalerna
      1 rotknöl
      1 rotknölar
      1 rotknölarna
      1 rotning
      2 rötning
      1 rötningen
      1 rots
      1 rotsaker
      1 rotstam
     18 rött
     25 rötter
      3 rotterdam
     14 rötterna
      1 rotundifolius
      1 rotytor
      1 rotz
      4 rouge
      1 roulette
      1 roulettehjul
      4 roundup
      1 roussimoff
      2 rouy
     14 rovdjur
      2 rovdjuren
      1 rovdjursbeteende
      1 rovfågels
      2 rovfåglar
      1 rovlevande
      1 rovor
      1 rövskrapor
      1 rowlings
      7 royal
      1 roz
      1 rozen
      1 rpk
      1 rpv
      1 rr
      1 rrintervall
      1 rrtid
      1 rs�[bensylpiperidylmetyl]dimetoxidihydroindenon
      1 rsc
      1 rsdioxopiperidinylhisoindolhdion
      1 [rshydroxioxofenylbutylhbensopyranon]
      1 rsmh
      1 rsmhrösträtt
      4 rsv
      4 rsvvirus
      3 rt
      1 rthämmare
      1 rtkorten
      4 rubbad
      1 rubbade
      2 rubbar
      1 rubbas
     17 rubbning
     16 rubbningar
      3 rubbningen
      4 rubella
      1 ruben
      2 rubens
      1 ruber
      1 rubescens
      1 rubinsteintaybis
      1 rubor
      2 rubra
      1 rubriceringar
      1 rubrik
      3 rubriken
      4 rubriker
      1 rubrikerna
      2 rubrum
      1 ruderatmarker
      1 rudi
      1 rüdiger
      1 rudiment
      1 rudimentär
      2 rudimentära
      9 rudolf
      1 ruess
      1 rugby
      1 rugbyspelare
      1 ruggat
      1 ruggig
      1 ruh
      2 ruiner
      1 ruinerad
      1 rule
      3 rulla
      1 rullade
      3 rullades
      2 rullande
      9 rullar
      2 rullarna
      6 rullas
      2 rullator
      2 rullats
      4 rulle
      1 rullen
      1 rullpapper
      1 rullstolen
     59 rum
      1 rumänen
      3 rumänien
      1 rumänsk
      1 rumänska
      1 rumbaprojektet
      1 rumens
      1 ruminanterbr
     11 rummet
      2 rummets
      2 rumsakustik
      1 rumsakustikern
      1 rumsdimensioner
      1 rumskamrater
      1 rumslig
      1 rumsligen
     18 rumstemperatur
      1 rumstempratur
      1 rumsväxt
      2 run
      1 runa
      1 runberg
      9 rund
     19 runda
     10 rundad
      5 rundade
      2 rundare
      1 rundat
      2 rundgång
      1 rundgått
      1 rundmask
     13 rundmaskar
      5 rundmaskarna
      1 rundmaskars
      1 rundmasken
      2 rundmunnar
      1 rundning
      1 rundnosade
      1 rundradions
      2 runge
      1 rungufolket
    206 runt
      6 runtom
      2 runtomkring
      4 ruptur
      1 rupturerade
      1 rupturerat
      1 rural
      1 rurala
      4 rus
      3 rusar
      1 rusdryck
      1 ruselii
      1 rusen
      5 ruset
      2 rusets
      1 rusframkallande
      3 rush
      2 ruska
      1 ruskan
      1 rusningstrafik
      1 russ
      1 russel
      3 russula
      1 russulaceae
      1 russyfte
      1 rusticus
      1 rustning
      1 ruston
      3 ruta
      2 rutan
      2 rutavdrag
      2 rutavdraget
      1 ruter
      3 ruterformad
      3 ruterformade
      1 ruterformen
      1 rutgersuniversitetet
      3 rutin
      1 rutinekg
      1 rutinen
     11 rutiner
      3 rutinerna
      2 rutinkontroll
      1 rutinkontrollen
      4 rutinmässig
      5 rutinmässiga
     13 rutinmässigt
      1 rutinsysselsättning
      2 rutinundersökning
      1 rutinvaccination
      3 rutmönster
      3 rutnät
      3 rutor
      1 rutten
      1 rutter
      1 ruttet
      1 ruttna
      1 ruttnande
      3 ruttnar
      1 ruttnat
      3 ruva
      1 ruvades
      2 ruvar
      2 ruvas
      1 ruy
      3 rv
      4 rvågen
      1 rvågens
      1 rvågor
      1 rw
      1 rwanda
      1 rxtechnology
      1 ryans
      1 ryck
      4 rycka
      1 ryckande
      6 rycker
      7 ryckiga
      6 ryckningar
      1 rycks
     24 rygg
      1 ryggar
      5 ryggbedövning
      5 ryggbesvär
      1 ryggbräda
     36 ryggen
      2 ryggens
      1 ryggkirurger
      2 ryggkirurgi
      4 ryggkotor
      3 ryggkotorna
      6 ryggläge
      1 rygglinje
      9 ryggmärg
     37 ryggmärgen
      3 ryggmärgens
      1 ryggmärgsbedövning
     12 ryggmärgsbråck
      1 ryggmärgsbråcksfall
      1 ryggmärgshinnorna
      1 ryggmärgskanalen
      1 ryggmärgsnerverna
      1 ryggmärgsprov
      1 ryggmärgssegment
      5 ryggmärgsskada
      1 ryggmärgsskador
      1 ryggmärgsstimulering
      7 ryggmärgsvätska
      4 ryggmärgsvätskan
      1 ryggmärgsvävnaden
      1 ryggmuskler
      2 ryggmusklerna
      1 ryggont
      1 ryggpartiet
      1 ryggproblem
      4 ryggrad
     36 ryggraden
      4 ryggradens
     21 ryggradsdjur
      3 ryggradsdjuren
      3 ryggradsdjurens
      1 ryggradsdjurs
     10 ryggradslösa
      1 ryggradsmanipulation
      1 ryggradssjukdomar
      1 ryggradsskada
      1 ryggradsskadade
      2 ryggsäck
      7 ryggskott
      1 ryggslutet
      6 ryggsmärta
      6 ryggsmärtor
      2 ryggsträng
      1 ryggsträngen
      1 ryggsträngs
      1 ryggsträngsdjur
      2 ryggvärk
      1 ryis
      9 rykte
      2 rykten
      3 ryktet
      1 rymd
      1 rymden
      1 rymdfarkoster
      1 rymdliftarkulturen
      1 rymdpromenader
      1 rymdresor
      1 rymdsjuka
      1 rymdsonder
      1 rymma
      1 rymmas
      6 rymmer
      1 ryms
      2 rymt
      1 rynkig
      7 rynkor
      1 rysk
      6 ryska
      4 ryske
      1 rysning
      1 rysningar
      2 ryssjukan
     28 ryssland
      9 rytm
      6 rytmer
      1 rytmgivare
      3 rytmisk
      4 rytmiska
      3 rytmiskt
      3 rytmrubbningar
      2 rytmstörningar
      1 ryttare
      1 ryttarens
      1 rzh�n
     43 s
      1 [s]
      4 sa
   2074 så
      1 saa
      1 saba
      1 sabbatsbergs
      1 sabelskenben
      1 saber
      1 sabina
      1 sabos
      1 sacer
      1 sachsska
      6 säck
      1 sackar
      1 sackarid
      3 sackarider
      1 sackarin
      1 sackaros
      1 säckig
      1 säcklik
      1 säcklika
      1 säckliknande
      1 säckmaskar
      1 saco
      1 sacroplasmisk
     10 säd
      1 sädadditiv
    143 sådan
    219 sådana
      1 sådande
     68 sådant
      1 sådd
      7 sade
      1 sadeh
      1 sadelnäsa
      6 säden
      3 sades
      1 sädesblåsa
      1 sädesblåsan
      1 sädesblåsesekret
      1 sädesblåsesekretet
      2 sädesblåsor
      2 sädesblåsorna
      4 sädesblåsornas
      1 sädescell
      1 sädescellen
      1 sädesceller
      1 sädesflytning
      1 sädesgrödor
      1 sädeskanaler
      2 sädeskanalerna
      2 sädesledare
      3 sädesledaren
      4 sädesledarna
      5 sädesslag
      1 sädesslagen
      1 sädessorter
      4 sädessträngarna
      3 sädesuttömning
      1 sädesuttömningar
     13 sädesvätska
      6 sädesvätskan
      1 sadistiska
      1 sadistiskt
      1 sadlar
      1 sadomasochism
      1 safarzadeh
      1 safavidiska
      1 safe
      1 saffires
      7 saft
      4 saften
      2 saftiga
      1 sag
     26 såg
      1 såga
    340 säga
      1 sågade
      1 sågades
      1 sagalitteraturen
      1 sagan
     23 sägas
      1 sagda
     48 säger
      2 sägnen
      1 sågning
      1 sågningen
      1 sagolik
      1 sågränna
     10 sågs
     52 sägs
     14 sagt
      3 sågtandad
      1 sågtandade
      1 sågtänder
      1 sågtandsmönster
      2 sagts
      3 sahachiro
      2 såhär
      7 sahara
      1 sahasrara
      8 sahlgrenska
      2 saint
      1 saintdizier
      1 saintlégerdepeyre
      1 saintlouis
      1 sainttropez
      1 sajter
     22 sak
      1 sakavdelningar
      4 saken
     81 saker
     36 säker
     32 säkerhet
      9 säkerheten
      3 säkerhets
      1 säkerhetsagenten
      1 säkerhetsarbete
      1 säkerhetsaspekter
      1 säkerhetsåtgärd
      1 säkerhetsåtgärder
      1 säkerhetsbedömning
      1 säkerhetsbetänkligheter
      1 säkerhetsbrister
      7 säkerhetsdatablad
      4 säkerhetsdatabladet
      1 säkerhetsexpertis
      1 säkerhetsfunktion
      1 säkerhetsgräns
      1 säkerhetsinformation
      1 säkerhetsklass
      1 säkerhetsklasser
      1 säkerhetskraven
      1 säkerhetsmärkningen
      2 säkerhetsmått
      1 säkerhetsmåttet
      1 säkerhetsnivån
      1 säkerhetsorgan
      1 säkerhetspolis
      3 säkerhetspolisen
      3 säkerhetspolitik
      1 säkerhetsregler
      2 säkerhetsrisk
      1 säkerhetsrisken
      1 säkerhetsrisker
      1 säkerhetsskäl
      1 säkerhetstester
      1 säkerhetstjänst
      2 säkerhetstjänster
      1 säkerhetsuppföljningen
      1 säkerhetsutbildningar
      1 säkerhetsutrustning
      1 säkerligen
      3 sakerna
     21 säkerställa
      2 säkerställas
      3 säkerställd
      2 säkerställda
      2 säkerställt
     49 säkert
      2 sakkunnig
      1 sakkunskap
      1 saklig
      7 sakna
      3 saknad
     13 saknade
      4 saknades
    114 saknar
     86 saknas
      2 saknat
     25 säkra
     12 säkrare
      1 säkras
      3 säkraste
      1 säkring
      1 sakroiliakaleden
      1 sakroilikalederna
      1 sakroplasmisk
     10 sakta
      3 saktar
      1 saktare
      1 sala
      2 salamander
      1 salamanderfamiljen
      1 salami
      1 sålänge
      5 sälar
      1 salbutamol
      1 salbutamolalbuterol
      5 sålda
      4 sålde
      1 såldedes
     22 såldes
      2 säldöd
      1 saldon
     68 således
      1 salem
      3 salen
      1 sälen
      2 salerno
      1 sälg
      1 salicylater
      1 salicylpreparaten
     10 salicylsyra
      1 salisb
     40 saliv
      2 salivavsöndring
      1 salivbrist
      1 salivdroppar
      8 saliven
      1 salivens
      1 saliveringen
      1 salivkörtlar
      1 salivutsöndring
      1 salix
     14 sälja
      1 säljare
      3 säljaren
     11 säljas
      7 säljer
     38 säljs
      1 sålla
      2 sallad
      1 sallader
      1 salladslök
    131 sällan
      1 sållar
      1 sållningsundersökningar
      5 sällskap
      3 sällskapet
      1 sällskaplighet
      7 sällskapsdjur
      1 sällskapsförening
     56 sällsynt
     69 sällsynta
      1 sällsyntare
      1 salmeterol
      2 salmiak
     12 salmonella
      1 salmonellaarter
      1 salmonellabakterier
      1 salmonellaepidemin
      1 salmonellainfektioner
      1 salmonellan
      1 salomon
      1 salomonöarna
      1 salongen
      2 salonger
      1 salpeteroxid
      8 salpetersyra
      1 salpetersyrans
      1 salpetersyrlighet
      1 salpingit
      1 salsa
      1 salsasåser
     47 salt
      3 sålt
      1 salta
      1 saltaktig
      2 saltartad
      1 saltbalansen
      1 saltbildning
      6 saltbrist
     26 salter
     15 saltet
      1 saltets
      1 saltfyndigheter
      2 saltgruvor
      3 salthalt
      1 salthaltig
      1 saltintaget
      1 saltkällor
      1 saltkristall
      1 saltkristaller
      1 saltlake
      1 saltlaken
      6 saltlösning
      1 saltlösningar
      1 saltrika
      5 sålts
      2 saltsug
     21 saltsyra
      4 saltsyran
      1 saltsyraproduktionen
      1 saltsyrasekretionen
      1 saltsyratillsats
      1 saltterapi
      8 saltvatten
      1 saltvattnet
      1 salubrin
      1 saluföra
      1 saluföras
      1 saluförda
      1 saluförde
      1 salufördes
      2 saluförs
      1 salufört
     15 sålunda
      2 salus
     10 salutogena
      6 salutogenes
     10 salva
      1 salvador
      1 salvadorii
      3 salvan
      1 salvare
     11 salvarsan
      1 salvarsanbehandlingarna
      1 salvarsanet
      1 salvarsanpreparatet
      1 salvform
      2 salvia
      9 salvor
      1 salzburg
      3 sam
      4 samarbeta
      6 samarbetade
      5 samarbetar
     27 samarbete
      5 samarbetet
      1 samarbetsmöjligheter
      1 samarbetsorganisationerna
      1 samarbetsproblem
      1 samarbetsprojekt
      1 samarbetsvillig
      1 samarium
      1 samart
      1 samba
    328 samband
      6 sambanden
     26 sambandet
      1 sambandstjänst
      1 sambladiga
      1 sambladigt
      2 sambuci
      1 sambucus
      2 sambunigrin
      2 sambyggare
      3 samer
      1 samernas
      2 sameskolan
      1 samevolution
      1 samexistera
      1 samexisterar
      1 samförekommer
      1 samförstånd
      1 samförståndet
      2 samfund
      1 samfunden
      1 samfundet
      1 samgraha
     25 samhälle
      6 samhälleliga
     23 samhällen
      1 samhällena
     78 samhället
     16 samhällets
      2 samhälls
      1 samhällsdiagnos
      1 samhällsekonomi
      2 samhällsfarliga
      6 samhällsförvärvad
      1 samhällsförvärvadaspiration
      1 samhällsförvärvade
      1 samhällsgemenskapen
      3 samhällsgrupper
      1 samhällsinstitution
      1 samhällsinstitutioner
      1 samhällsklasserna
      1 samhällskostnad
      1 samhällskostnaderna
      1 samhällsmakten
      2 samhällsmedicin
      1 samhällsmoral
      2 samhällsnivå
      1 samhällsordning
      1 samhällsperspektiv
      2 samhällsplanering
      1 samhällspreventiv
      1 samhällsstress
      1 samhällsstrukturen
      1 samhällsstrukturens
      1 samhällsstrukturer
      1 samhällssynen
      1 samhällssystemet
      1 samhällsvetenskapen
      2 samhällsvetenskapliga
      4 samhita
      1 samhitas
      2 samhörande
      3 samhörighet
      3 saminfektion
      1 saminofenylpropanon
      1 samiskans
      1 samkhya
      1 samkhyatraditionen
      2 samklang
      4 samkönade
     14 samla
      3 samlad
     13 samlade
      1 samlades
     90 samlag
      2 samlagen
      5 samlaget
      1 samlagsexuella
      1 samlagssmärtor
      2 samlagsställningar
      3 samlande
     14 samlar
      4 samlare
      1 samlarfolk
      1 samlarföremål
      1 samlarsamhällen
      1 samlarvärdet
     27 samlas
      1 samläser
      2 samlat
      7 samlats
      1 samlevnad
      1 samlevnadsundervisning
     13 samling
      1 samlingar
      1 samlingbeteckning
      5 samlingsbegrepp
      1 samlingsbenämning
      2 samlingsbeteckning
      2 samlingskondom
     40 samlingsnamn
      4 samlingsnamnet
      1 samlingsordet
      1 samlingsplats
      1 samlingsrör
      1 samlingswebbplatsen
      1 samliv
      1 samlivet
    470 samma
     84 samman
      1 sammanband
      1 sammanbinda
      1 sammanbinder
      1 sammanblanda
      3 sammanblandas
      1 sammanbunden
      2 sammanbundna
      5 sammandragande
      1 sammandraget
      2 sammandragna
      7 sammandragning
      6 sammandragningar
      1 sammandragningarna
      3 sammandragningen
      1 sammandras
      1 sammanfall
      1 sammanfalla
      3 sammanfallande
      8 sammanfaller
      3 sammanfattade
      1 sammanfattades
      6 sammanfattande
      3 sammanfattar
      1 sammanfattas
      2 sammanfattat
      2 sammanfattning
      1 sammanfattningen
      2 sammanfattningsvis
      1 sammanflätade
      1 sammanflöde
      2 sammanfoga
      1 sammanfogade
      1 sammanfogar
      3 sammanfogas
      1 sammanfogningar
      1 sammanfogningarna
      1 sammanförda
      2 sammanförs
      1 sammanhållande
      2 sammanhållna
      1 sammanhållningen
      1 sammanhålls
    102 sammanhang
      8 sammanhängande
      1 sammanhangen
     19 sammanhanget
      1 sammankokade
      1 sammankoppla
      2 sammankopplad
      2 sammankopplade
      1 sammankopplar
      1 sammankopplas
      3 sammankopplat
      2 sammankopplats
      3 sammankoppling
      2 sammankopplingen
      1 sammanlagd
      3 sammanlagda
      1 sammanlagras
      2 sammanlagringsfri
     12 sammanlagt
      1 sammanlänkad
      3 sammanlänkade
      1 sammanlänkas
      1 sammanliknar
      7 sammansatt
     11 sammansatta
     24 sammansättning
      1 sammansättningaktivitet
      2 sammansättningar
      4 sammansättningen
      1 sammanslagen
      3 sammanslagning
      1 sammanslagningen
      2 sammansmälta
      1 sammansmälter
      2 sammansmältning
      2 sammansmältningen
      4 sammanställa
      1 sammanställas
      1 sammanställd
      1 sammanställda
      3 sammanställdes
      4 sammanställer
      5 sammanställning
      1 sammanställningen
      4 sammanställs
      2 sammanställt
      1 sammantagen
      9 sammantaget
      3 sammantagna
      1 sammanträden
      2 sammanträder
      1 sammanträffande
      1 sammantryckta
      1 sammanvägning
      3 sammanväxningar
      1 sammanväxningaradherenser
      1 sammanväxta
      1 sammanviga
      3 sammanvuxna
      2 samme
      1 sammet
      1 sammetsblomster
      1 sammetssvart
      1 sammoniak
      2 samordna
      2 samordnande
      2 samordnar
      1 samordnas
      1 samordnat
      1 samordnats
      3 samordningsansvar
      2 samordningsansvaret
      1 samordningsgrupp
      1 samp
      1 samplar
      1 samples
      1 sampling
      1 samplingsfrekvensen
      1 sampolymer
      7 samråd
     50 sämre
      2 samröre
      2 samsara
      9 samsjuklighet
      1 samsö
     23 samspel
      2 samspela
      1 samspelar
      8 samspelet
      1 samspelets
      1 samspelkommunikation
      1 samspelsmönstret
      1 sämst
      4 sämsta
      1 samstämmiga
      2 samstämmighet
      1 samstämmigheten
      4 samsyn
    869 samt
     19 samtal
      4 samtala
      4 samtalen
      3 samtalet
      1 samtals
      9 samtalsterapi
      1 samtalsterapin
      1 samtid
      9 samtida
      1 samtiden
      1 samtidens
     13 samtidig
      4 samtidiga
    173 samtidigt
     80 samtliga
      2 samtyckande
      9 samtycke
      1 samtycker
      1 samtyckesdokument
      1 samtyckt
      7 samuel
      1 samuelsgatan
      2 samurajer
      1 samvariation
      1 samvariera
      3 samvaro
      3 samverka
     18 samverkan
      1 samverkande
      1 samverkansarbetet
     17 samverkar
      3 samvete
      1 samvetsgrant
      1 samvetsömhet
      2 san
      1 sanatoriebyggnaden
      1 sanatoriekuren
      1 sanatorieläkare
      2 sanatoriemiljön
     11 sanatorier
      6 sanatorierna
      5 sanatoriet
      1 sanatoriets
      1 sanatorievård
      6 sanatorium
      1 sanct
      1 sancti
      3 sand
      4 sända
      4 sändare
      1 sändarspole
      1 sandberg
      1 sandblästring
      1 sande
      1 sände
      2 sändebud
      1 sandell
      1 sandemos
      2 sanden
     18 sänder
      5 sändes
      1 sandfång
      1 sandfånget
      1 sandfärgadbeige
      1 sandfilter
      1 sandfly
      2 sandig
      1 sandiga
      1 sandin
      2 sandjord
      1 sandkorn
      1 sandlåda
      1 sandlådesjukan
      1 sandmyggefeber
      2 sandmyggor
      1 sändning
      1 sandoz
      3 sandpapper
      1 sandpappersfilar
     12 sänds
      1 sandstormar
      1 sandstranden
      1 sandstränder
      1 sandträsk
      1 sandvikens
      1 sandwicensis
      1 sane
      2 sanerar
      1 sanerare
      1 saneraren
      2 saneras
      6 sanering
      1 saneringrivningborttagande
      3 saneringsbolag
      1 sanfranciscensis
     12 sång
      1 säng
      2 sängar
      1 sångare
      1 sängbäcken
      1 sängbenen
      1 sängbord
      1 sängbunden
      1 sängbundna
      1 sängelag
      1 sången
     19 sängen
      2 sanger
      1 sänger
      2 sångerskan
      1 sängkamrater
      1 sängkanten
      6 sängkläder
      5 sängläge
      4 sängliggande
      1 sångmikrofon
      3 sängrökning
      3 sängs
      1 sångsammanhang
      1 sångteknik
      2 sanguinaria
      1 sanguinolentum
      1 sängvätande
      4 sängvätare
     11 sängvätning
      1 sängvätningen
      1 sangviniskt
      1 sangvinska
      1 sanhansurta
      2 sanitaire
      1 sanitära
      1 sanitation
      5 sanitet
      2 sanitetsåret
      1 sanitetsområden
      1 sanitetssystem
      1 sanitetsvaror
      1 sanitoriekomplexen
      1 sanity
      1 sank
     32 sänka
      7 sänkan
      1 sänkas
      1 sänkbara
      2 sanke
     28 sänker
      8 sänkning
      1 sänkningen
      2 sänkningsreaktion
      1 sänkningsreaktionen
      1 sänkningsreaktionens
      1 sänkningsvärdet
      7 sänks
      3 sankt
     28 sänkt
     14 sänkta
      1 sänkte
      1 sänktes
      1 sanktioner
      1 sanktionerade
      1 sanktionerades
      1 sänktmedvetandegrad
      1 sann
      8 sanna
      2 sanning
      1 sanningar
      3 sanningen
      1 sanningsanspråk
      1 sanningsdrog
      1 sanningsenliga
      2 sanningsserum
      3 sannolik
      3 sannolikast
     17 sannolikhet
     31 sannolikheten
      1 sannolikhetsskala
     58 sannolikt
      1 sano
      1 sanofi
      1 sans
     11 sanskrit
      1 sanskritord
      2 sanskritordet
      1 sanskrits
      4 sant
      1 santa
      1 santarelli
      1 santiago
      1 santonin
      1 santoriefrågan
      1 saob
      4 såpa
      2 såpass
      1 säper
      1 sapfoe
      1 sapiens
      1 såplösning
      1 såplut
      1 såpnejlika
      1 såpnejlikan
      1 saponaria
      1 saponifiering
      1 saponiner
      1 säpos
      1 sapotace�
      1 sapotaceae
      1 sapovirus
      1 saprofyticus
      1 saprophyticus
      1 saptadhatu
     63 sår
      1 såra
      1 sårad
      6 sårade
      1 säras
      1 sarasdjinjasstammen
      1 saraswati
      1 sårat
      1 sårbakterier
      1 sårbar
      2 sårbara
      1 sårbarare
      6 sårbarhet
      3 sårbarheten
      1 sårbarheter
     11 sårbarhetsmodellen
      4 sårbehandling
      1 särbehandling
      2 sårbildning
      1 sårbotten
      2 sarcom
      2 sarcos
      1 sårdesinfektion
      1 sardinien
      1 sardonicus
      1 särdrag
      1 särdragen
      1 särdraget
      1 säregna
      8 såren
     35 såret
      2 sårets
      1 sårfebrar
      2 sårig
      2 såriga
     12 sarin
      1 sarinångor
      1 sarinattack
      1 sårinfektioner
      2 sarinförgiftning
      1 saringas
      1 saringasattacken
      1 saringasen
      1 sark
      2 sårkanterna
      4 särklass
      7 sarkoidos
      1 sarkoidosen
      1 sarkoidossom
     22 sarkom
      1 sarkomassocierat
      1 sarkomvarianten
      1 sarkopeni
      6 sårläkning
      1 sårnader
      1 sarno
      1 sårodling
      1 sårpenetrerande
      1 särpräglade
      8 sars
      1 sårsjukdomar
      2 sårskada
      1 sårskadan
      3 sårskador
     70 särskild
     66 särskilda
     14 särskilja
      1 särskiljandet
      2 särskiljas
      5 särskiljer
      1 särskiljs
    300 särskilt
      2 särskola
      3 särskolan
      1 särskolans
      2 särskoleelever
      1 särskoleläkaren
      1 sårskorpor
      1 särskrivning
      1 sårtejp
      1 sårtvätt
      1 sårvård
      1 sårvätska
      1 sårvätskor
      1 sårvävnad
      2 sarvimäki
      1 särvux
      1 sås
      1 sasaniderna
      1 [sasch]
      1 såser
      2 sashimi
    401 såsom
      1 såsomnaegleria
      4 säsong
      1 säsongbunden
      1 säsongen
      1 säsongs
      1 säsongsbetonade
      1 säsongsbunden
      1 säsongsgrönsaker
      1 sastrawan
      1 satanas
      1 satans
      2 satchidananda
      1 satdaghensis
      6 säte
      1 satellitstater
      1 satellitteknologi
      2 säters
      2 sätesbjudning
      1 sätesmuskler
      1 sätet
      1 såtillvida
      1 satir
      1 satiriska
      1 sativa
      1 sats
      3 satsa
      1 satsade
      3 satsar
      1 satsas
      1 satsat
      1 satsbyggnad
      1 satsmelodi
      1 satsning
      1 satsningar
      1 satsningen
      1 satstestning
     23 satt
    535 sätt
      1 satta
     39 sätta
     24 sättas
      8 satte
      6 sätten
     37 sätter
      8 sattes
     43 sättet
      1 sättningar
      1 sättpotatis
      7 satts
     77 sätts
      1 saturated
      1 saturationen
      1 saturationsmätare
      1 saturnism
      1 saturnus
      3 saudiarabien
      1 sauer
      1 saul
      3 sauna
      1 saunominen
      2 saureus
      1 sauternesviner
      1 sav
    122 såväl
      1 savanner
      1 savant
      5 sävenbom
      1 sävenbomolja
      1 savi
      2 såvida
      2 såvitt
      1 sävsjö
      1 savusauna
      1 saxatilis
      1 saxliknande
      1 saxofonisten
      3 saxon
     21 sbu
      2 sca
      1 scaevola
      2 scala
      1 scalaris
     11 scale
      1 scan
      1 scandinavian
      1 scannar
      1 scarlett
      1 scb
      1 scbs
      2 sceller
      2 scen
      1 scenario
      2 scenen
      1 scener
      1 scenframträdanden
      5 scenkonst
      1 scenkonstnärinna
      1 scenskräck
      2 scf
      1 schaarschmidt
      2 schack
      1 schackspel
      3 schäfer
      1 schäfrar
      2 schaktugnar
      7 schaman
      9 schamanen
      4 schamaner
      2 schamanerna
      1 schamaniska
      5 schamanism
     12 schamanismen
      1 schamanismens
      4 schamanistiska
      1 schamans
      1 schamanska
      1 schamanskt
     12 schampo
      4 schampon
      1 schamponeringsmedel
      1 schamposorter
      2 schampot
      4 schanker
      2 schankern
      1 schappel
      1 scharlakansbär
      3 scharlakansfeber
      2 schaudinn
      1 schaumanns
      1 schedule
      1 scheele
      3 scheibel
      1 scheibels
      1 schellhas
      4 schema
      1 schemalagda
      1 schemalägga
      2 schemat
      1 schematisk
      1 schematiskt
      1 scheppel
      1 schimpans
      4 schimpanser
      1 schimpanskadaver
      1 schinz
      1 schismer
      1 schismerna
      4 schistosoma
      7 schistosomiasis
      1 schitzofrena
      2 schizo
      2 schizoaffektivt
      2 schizofren
     13 schizofrena
    255 schizofreni
      2 schizofrenia
      5 schizofrenidiagnos
      2 schizofrenidiagnosen
      2 schizofrenidiagnoser
      1 schizofrenidiagnostiken
      1 schizofrenidiagnostisering
      1 schizofreniepisoder
      2 schizofrenier
      3 schizofrenierna
      8 schizofreniliknande
      4 schizofrenin
      1 schizofrenins
      1 schizofrenis
      1 schizofrent
      2 schizont
      1 schizonten
      1 schizonter
      1 schizonterna
      1 schizosaccharomyces
      1 schizotyp
      1 schizotypa
      1 schizotypi
      2 schlesien
      1 schnalstal
      1 schneibel
      1 schneider
      1 schoenbuchensis
      1 schönbein
      1 schöningen
      1 schöningerspjuten
      1 schönlein
      5 school
      5 schopenhauer
      1 schrader
      1 schrothmetoden
      1 schubert
      1 schuur
      1 schwabiska
      1 schwannska
      8 schweiz
      2 schweizaren
      2 schweizisk
      4 schweiziska
      2 schweiziske
      1 schyman
     18 science
      1 sciencefictionartade
      5 sciences
      1 scientific
      2 scintigrafi
      1 scintillation
      1 scintillationseffektivitet
      2 scintillatorer
      1 sclera
      1 scombroidförgiftningen
      1 scombroidosis
      1 scopolia
      4 score
      2 scoring
      3 scott
      1 scouter
      1 scouternas
      1 scq
      3 scrapie
      1 scream
      6 screena
      1 screenades
     15 screening
      1 screeningapparaten
      1 screeninghänseende
      6 screeningprogram
      1 screeningprogrammet
      1 screeningsmetoder
      1 screeningtest
      1 screeningtester
      1 screeningundersökning
      1 screeningundersökningar
      1 scrooge
      1 scrotum
      2 scs
      1 sct
      1 scuman
      1 scutellatus
      2 sd
      1 sda
      1 sdb
      1 sdelen
    385 se
      1 seal
      1 seattle
      2 sebastian
      1 sebek
      2 seborré
      1 seborrhoeic
      4 seborroisk
      1 seborroiska
      3 seborroiskt
      1 sebum
      2 secale
      1 secaliner
      1 secam
      2 second
      2 secondhandföremål
      1 secondhandmöbler
      1 secret
      2 sectio
      1 securitas
      2 sécurité
      1 security
      5 sed
    737 sedan
      2 sedativ
      2 sedativa
      1 sedativum
      2 sedda
      1 sedens
      1 seder
      2 sederande
      5 sedering
     17 sedermera
      1 sederna
      1 sedesfördärv
      1 sedgwick
      1 sedibus
      1 sediment
      1 sedimentation
      1 sedimentationsbassäng
      1 sedimentera
      1 sedimenterar
      1 sedimenteras
      2 sedimentering
      1 sedimenteringen
      2 sedimenteringsbassängen
      1 sedimenteringsförtjockaren
      2 sedimenteringsproblem
      1 sedlar
      1 sedmintationshastoghete
      1 sednan
      2 sedvänjan
      3 sedvanlig
      1 seelenkunde
      6 seende
      1 seendet
      1 seendets
      1 seg
      1 sega
      3 segel
      1 segelklaffarna
      1 segelsättning
      1 seger
      1 segerhuva
      1 seglande
      1 seglar
      1 seglats
      2 seglet
      9 segment
      1 segmentduration
      2 segmenten
      1 segmentera
      3 segmenterade
      1 segmenteras
      1 segmentering
      1 segmenteringen
      1 segmentet
      1 segraren
      1 segré
      1 segregering
      7 segt
      1 segue
     13 segway
      1 segways
      1 seitan
      1 sej
      1 sejd
      1 sejdat
      1 sejin
      1 sek
      1 sekalin
      1 sekel
      5 sekelskiftet
      1 sekelvända
      1 sekentei
      2 sekler
      2 seklet
      1 sekonden
     27 sekret
      2 sekretesskyddet
      1 sekretets
      8 sekretin
      1 sekretinet
      6 sekretion
      1 sekretionen
      2 sekretorisk
      1 sekretoriska
      2 sekt
      3 sekten
      1 sektens
      1 sekter
      5 sektion
      2 sektionen
      2 sektionnätverk
      1 sektliknande
      3 sektor
      1 sektorer
      1 sektoriell
      3 sektorn
      1 sekulär
      1 sekulariserade
     12 sekund
     47 sekundär
     43 sekundära
      1 sekundärcancer
      1 sekundärfall
      1 sekundärfolliklarna
      2 sekundärgranula
      1 sekundärinfekterade
      1 sekundärinfekteras
      1 sekundärinfektion
      1 sekundärprevention
      1 sekundärsmitta
      1 sekundärstadiet
      1 sekundärstruktur
     11 sekundärt
      2 sekunden
     21 sekunder
      1 sekunder�
      1 sekunderna
      1 sekunderruta
      1 sekundsnabba
      2 sekvens
      3 sekvensen
      2 sekvenser
      3 sekvensering
      1 sekventiellt
      1 selarbetet
      1 seldinger
      1 seldingerteknik
      3 sele
      1 selection
      3 selegilin
      1 selegilinet
      1 selekteras
      2 selektion
     11 selektiv
     11 selektiva
      2 selektivitet
      1 selektivitetsfilter
      1 selektivt
      4 selen
      1 selfdefeating
      1 selfinjury
      2 seligman
      2 seligmans
      2 selikoff
      2 sella
      1 selleri
      1 selleripersilja
      2 selman
      1 selye
      1 semantik
      1 semantisk
      1 semenis
      1 semester
      1 semesteranläggningar
      6 semg
      1 seminandi
      2 seminarier
      1 seminiferous
      1 seminom
      2 semipermeabelt
      1 semistrukturerad
      1 semitransparent
      3 semivegetarianer
      1 semmelweis
      4 semmelweiss
      1 sempers
     47 sen
     18 sena
      2 senan
      1 senans
      1 senap
    454 senare
      1 senares
     14 senast
     74 senaste
      1 sendebuterande
      1 sendoxan
      1 seneca
      2 senegal
      1 senescens
      2 senfästen
      1 senfästesinflammation
      1 senfästesinflammationerna
      1 senförflyttningar
      1 senförlängningar
      2 senhet
      3 senil
      2 senildemens
      1 senilis
      2 senilitet
      2 seniorboende
      1 seniorboendettrygghetsboendet
      1 senis
      1 senlatin
      1 senlatinets
      1 senmedeltiden
      1 senna
      5 senor
      1 senreflexer
      1 senrenässansen
      1 sens
      1 sensationen
      2 sensationer
      2 sense
      1 senseartat
      2 sensibiliserad
      1 sensibiliserande
      1 sensibilitetsnedsättning
      1 sensitiseras
      2 sensitisering
      1 sensitiseringen
      1 sensitiv
      1 sensitiva
      2 sensitive
      9 sensitivitet
      2 sensitivity
      1 sensitivt
      1 sensivitet
      2 sensommaren
      2 sensomotoriska
      4 sensor
      1 sensoranalys
      1 sensorer
      1 sensorik
      1 sensorineural
     16 sensorisk
     30 sensoriska
      1 sensorisktmotoriskt
      1 sensoryseeking
      1 sensuell
     47 sent
      1 sentao
      3 sentida
      1 senvintern
      2 senytorna
      1 sep
      1 separarera
      8 separat
      9 separata
      1 separationen
      1 separationer
      4 separationsångest
      1 separationsmetod
      1 separationsprocess
      1 separationsteknik
      9 separera
      1 separerad
      2 separerade
      1 separerades
      6 separerar
      7 separeras
      2 separerat
      2 separerats
      1 sephadex
      1 seppuku
     41 sepsis
      1 sepsispatienter
     27 september
      1 septembermorden
      1 septentrionale
      2 septikemi
      5 septisk
      7 septum
      2 septumpiercing
      1 septumpiercingar
      2 septumpiercingen
      1 septumpiercingstraditioner
      1 sequence
    187 ser
      1 sera
      2 serafimerlasarettet
      1 serafimerordensgillet
      1 serafimerordenslasarettet
      1 serafimerriddare
      2 serdolect
      1 serge
      1 sergej
      1 sergey
      2 serial
     19 serie
      1 seriefigur
      1 seriefiguren
      1 seriekopplade
      1 seriemördare
      7 serien
      1 serienummer
      4 serier
      1 serierna
      2 serietidningar
      1 serietillverkade
      2 seriös
      3 seriösa
      1 serm
      4 serologi
      2 serologisk
      3 serologiska
      2 serologiskt
      1 seronegativa
      1 seropositiva
      1 serös
      1 serösa
      1 seröst
      1 serotonerg
      1 serotonerga
      2 serotonergt
     27 serotonin
      1 serotoninaktivitet
      1 serotoninåterupptagningshämmaren
      4 serotoninåterupptagshämmare
      1 serotoninbalans
      1 serotonindopaminbalansen
      1 serotoninets
      1 serotoninhalten
      1 serotoninhypotesen
      1 serotoninreseptorer
      1 serotoninsystem
      4 serotyp
      1 serotypen
      6 serotyper
      4 serotypspecifika
      1 seroxat
      2 serpentin
      1 serpentina
      1 serpyllifolia
      5 sertindol
      2 sertoliceller
      1 sertolileydigcellstumör
      1 sertralin
      1 serullas
     12 serum
      1 serumelektrolyter
      1 serumet
      1 serumglukos
      1 serumkreatinin
      1 serumvärden
      1 serva
      4 serveras
      1 servering
      1 serveringsställen
      1 servett
      1 servetten
     17 service
      1 servicebranschen
      1 servicebranschens
      1 servicehund
      1 servicehus
      1 serviceinsatser
      1 servicepersonal
      2 services
      1 servier
      1 serviser
      1 servitör
    159 ses
      1 sesam
      1 session
      1 sessionerna
      1 sestamibi
      1 set
      1 setifolius
    149 sett
      9 setts
      1 sevesokatastrofen
      3 sevofluran
      1 sevoflurane
    131 sex
      3 sexarbetare
      1 sexarbete
      1 sexårig
      1 sexberoende
      1 sexcentrum
      1 sexdagar
      1 sexistisk
      1 sexköpslagen
      1 sexlingar
      1 sexliv
      2 sexlust
      1 sexmånader
      1 sexobjekt
      1 sextalig
      1 sexterapeut
      1 sexterapi
      1 sextio
      1 sextiotal
      1 sextiotalistgenerationen
      3 sexton
      1 sextondelar
      1 sexual
      5 sexualbrott
      1 sexualbrottsrubriceringarna
      2 sexualdriften
      1 sexualförbrytare
      1 sexualiserad
      9 sexualitet
      6 sexualiteten
      1 sexuallivet
      1 sexualmorals
      1 sexualpartnern
      1 sexualskräck
      1 sexualvaneundersökning
     66 sexuell
     58 sexuella
     63 sexuellt
      1 sfa
      2 sfär
      1 sfären
      1 sfärisk
      3 sfäriska
      1 sfäriskt
      1 sfe
      1 sfetibc
      1 sfinkter
      1 sfinktrarna
      1 sform
      1 sformad
      2 sformen
      1 sfrf
      4 sfs
      1 sfsr
      1 sgs
      1 sgu
      1 shadow
      1 shaiva
      1 shakerssekten
      1 shakesen
      1 shakespeare
      1 shakespeares
      1 shakti
      1 shaktiton
      1 shaman
      1 shamanen
      3 shamaner
      1 shamanerna
      1 shamaners
      1 shamanistiska
      1 shambhala
      1 shampooing
      1 shampots
      1 shang
      1 shanghai
      5 shangrila
      1 shankle
      2 shapiro
      1 sharia
      1 sharialagar
      1 sharp
      1 sharpeyschafer
      1 shatkarma
      1 shaw
      2 shawpriset
      1 shbam
      3 shbg
      1 shbgnivåerna
      1 sheanötter
      2 shearwave
      1 sheasmör
      4 sheasmöret
      1 sheasmörets
      1 shela
      2 shelby
      1 shell
      1 sheminvägen
      1 sheriff
      1 sheriffer
      1 sherlock
      4 shiatsu
      1 shiatsumassör
      1 shiatsutekniken
      1 shibasaburo
      1 shields
      2 shift
      1 shiga
      1 shigatoxin
      5 shigella
      1 shigellos
      1 shikimicsyra
      1 shimon
      1 shimpanser
      2 shin
      1 shiner
      1 shinrikyo
      1 shinto
      1 shintoismen
      1 shintōmytologi
      1 shirley
      2 shiva
      1 shmerlings
      4 shock
      1 shogunatet
      1 shoot
      1 shorts
      1 show
      1 shown
      1 shprintzen
      1 shprintzens
      1 shramanatraditionerna
      2 shrodes
      1 shudo
      1 shukra
      1 shumway
      6 shunt
      1 shuntas
      1 siadh
      1 sialinsyra
      1 siamesiska
      5 sibirien
      4 sibutramin
      4 sicilien
      3 sick
      1 sickel
      1 sickelcellanemi
      1 sickelcellsanemi
      4 sickle
      2 sicklecellanemi
      3 sickness
      1 si�clefatalism
      1 siculus
      6 sid
     68 sida
    100 sidan
      1 sidans
      3 sidas
      3 siden
      2 sidenbaner
      1 sidiplattan
      1 sidkedjan
      1 sidkrafter
      2 sidkrafterna
      4 sidled
      1 sidney
      1 sidnummer
      1 sidoaxlar
      1 sidobetydelse
      1 sidoeffekt
      3 sidoeffekter
      1 sidoeffekterna
      2 sidogren
      1 sidogrenarna
      1 sidogrupper
      1 sidokedja
      3 sidokedjor
     19 sidor
     15 sidorna
      1 sidorötter
      1 sidoskalmar
      1 sidoväggarna
      1 sidovapen
      2 sidvind
      1 siegel
      1 siegemundin
      1 siegmund
      1 siemerlingcreutzfeldt
      1 sienhet
      3 sienheten
      1 sienheter
      4 sierra
      5 sievers
     11 sievert
      1 sifferbeteckningen
      1 sifferfakta
      1 siffertecken
      1 siffertecknet
     15 siffra
     18 siffran
     14 siffror
      7 siffrorna
      3 sifneos
   2546 sig
      1 sigault
      1 sighsten
      1 sigill
      1 sigmoid
      1 sigmoidala
      2 sigmoideoskopi
     23 sigmund
     20 signal
      1 signalämne
      1 signalbearbetningen
      2 signalbehandling
      1 signaldetektering
     23 signalen
      2 signalens
     82 signaler
      1 signalera
      2 signalerande
     12 signalerar
      2 signalering
      1 signaleringen
     13 signalerna
      1 signalernas
      1 signalers
      1 signalförmedling
      1 signalfrekvensen
      1 signalgenerator
      1 signalgeneratorer
      1 signalmolekyl
      3 signalöverföring
      3 signalöverföringen
      1 signalproteinerså
      1 signalreaktion
      1 signalspektrumet
      7 signalsubstans
      4 signalsubstansen
     17 signalsubstanser
      2 signalsubstanserna
      1 signalsystem
      1 signalsystemet
      1 signaltransduktor
      2 signalupptagning
      3 signaturläran
      1 signe
      1 signerar
      1 signerier
      1 signetics
      2 signifikans
      1 signifikansen
      1 signifikansnivån
      1 signifikanstester
     23 signifikant
      1 sigrid
      1 sigur
      1 sik
     35 sikt
      1 siktande
      1 siktar
      1 sikten
      2 sildenafil
      1 silederna
      1 silene
      1 siler
      1 silhuett
      1 silhuetten
      1 siliconhydrogelmaterial
      1 silikat
      1 silikater
      2 silikatmineral
     10 silikon
      1 silikonbelagda
      1 silikonbelagdahydrogelbelagda
      1 silikonet
      1 silikonkateter
      1 silikonplatta
      1 silikonplattan
      1 silikonproteser
      1 silikonproteserna
      1 silikonskål
      8 silikos
      1 silikosknutor
      3 silke
      1 silkesfjärilen
      1 silkesglänsande
      1 silkesnäsdukar
      1 silmo
      4 silor
      1 silva
     16 silver
      1 silverbelagda
      1 silvereternell
      2 silverfärgad
      1 silverframställning
      3 silverframställningen
      1 silverglasögon
      1 silvergruva
      1 silvergruvorna
      1 silverhalid
      2 silverhalider
      1 silverhalidfällning
      4 silverjodid
      3 silverklorid
      1 silverkrut
      1 silvernät
      9 silvernitrat
      1 silveroxid
      1 silversalt
      1 silversalter
      1 silvertip
      2 silvervit
      1 silvervitt
      1 silvias
      1 silvrets
      1 sim
      1 simbassänger
      1 simförmåga
      2 simhallar
      1 simhopp
      1 simhud
      1 simila
      1 similar
      2 similia
      3 similibus
      6 simma
      1 simmande
      3 simmar
      1 simmarklåda
      7 simning
      4 simon
      1 simonfokus
      1 simopoulos]
      1 simövningen
      1 simpel
      4 simplex
      5 simplexvirus
      1 simplicity
      1 simponi
      1 simpson
      1 simri
      1 simrörelser
      1 simson
      1 simsträcka
      1 simtur
      1 simturer
      2 simulator
      4 simulera
      3 simulerad
      1 simulerade
      1 simulerat
      2 simulering
      1 simuleringsverktyg
      1 simulium
      1 simultan
    805 sin
    424 sina
      1 sinaftin
      1 sinaloa
      1 sindbisvirus
      1 sindh
      1 sine
      1 sinead
      1 sinéad
      3 sing
      2 singalerar
      5 singapore
      1 singel
      1 singer
      1 singh
      3 singular
      1 singularform
      1 singularis
      1 sinister
     10 sinne
      1 sinnelag
     13 sinnen
      7 sinnena
      1 sinnesapparater
      1 sinnesavvikelser
      1 sinnesceller
      3 sinnesförnimmelser
      1 sinneshåren
     27 sinnesintryck
      3 sinnesintrycken
      1 sinnesintrycket
      1 sinnesmodaliteterna
      1 sinnesnervbanor
      1 sinnesorgan
      2 sinnesorganen
      2 sinnesrörelse
      1 sinnessignaler
      1 sinnessjuka
      4 sinnessjukdom
      2 sinnessjukhus
      1 sinnessjukhusen
      1 sinnessjuklagstiftningen
      5 sinnesslö
      4 sinnesslöa
      2 sinnesslöhet
      5 sinnesstämning
      3 sinnesstämningar
      3 sinnesstämningen
      1 sinnesstimuli
      1 sinnessystem
      1 sinnestämningen
      2 sinnestillstånd
      1 sinnestillståndet
      1 sinnesundersökningar
      1 sinnesupplevelse
      1 sinnesupplevelsen
      5 sinnesupplevelser
      1 sinnesupplevelserna
      1 sinnesvillor
      4 sinnet
      1 sinnets
      3 sinsemellan
      1 sinuatum
      5 sinuit
      1 sinuitsinusit
      9 sinus
      2 sinusarrytmi
      1 sinusbesvär
      1 sinusbradykardi
      1 sinusformade
      1 sinusknuta
      7 sinusknutan
      1 sinuskurvor
      2 sinusoider
      6 sinusrytm
      3 sinusrytmen
      2 sinussyndrom
      1 sinustakykardi
      1 siotetraherar
      1 siphonaptera
      1 sippan
      2 sipporna
      2 sippra
      1 sipprar
      2 sippsläktet
      8 sir
      2 sirap
      1 sirapslösningar
      3 sirenomelia
      2 sirs
      1 sirsinfektion
      1 sis
      1 sisådär
      1 sisal
      1 sisalagave
      1 sisalana
      1 sisohsas
     10 sist
     58 sista
      2 siste
     21 sistnämnda
      1 sistnämnde
      1 sisu
      1 sisyfos
      1 sit
      1 site
      1 sites
      3 sits
    355 sitt
     37 sitta
     12 sittande
      1 sittandes
      4 sittbad
    137 sitter
      1 sitterligger
      2 sittning
      1 sittplats
      1 sittposition
      1 sittringen
      2 sittställning
     10 situ
     44 situation
      1 situationella
     27 situationen
     60 situationer
      1 situationerna
      1 situationsberoende
      1 situationsbetingad
      1 situaton
      1 situcancern
      1 siugdom
      1 sivananda
      1 sivlér
      1 six
      1 size
      1 sj
     34 själ
      1 själamässorna
      1 sjalar
      4 själar
      2 själarna
      1 själavandring
      1 själavård
     27 själen
      6 själens
      1 själland
      1 själlandskrönikan
      1 själpsyke
      4 själsbegreppet
      1 själsförmögenheterna
      3 själsliga
      1 själsligt
      2 själslivet
      1 själstillstånd
    248 själv
    228 själva
      1 självadministrering
      1 självalstrat
      1 självannan
      1 självantänder
      1 självbalanserande
      1 självbefruktas
      1 självbehandling
      1 självbehärskning
      2 självbestämmande
     16 självbild
      4 självbilden
      1 självbiografiskt
      1 självdestruktiva
      2 självdestruktivitet
      5 självdestruktivt
      1 självdialyspatienter
      1 självdisciplin
      1 självdråparen
      5 självet
      1 självfertila
      1 självförebråelse
      1 självförhärligande
      1 självförnyande
      1 självförsjunkenhet
      1 självförsörjande
      1 självförståelse
      1 självförsvar
      1 självförsvarsvapen
      4 självförtroende
      1 självförtroendet
      1 självförvållad
      1 självförvållade
      3 självförverkligande
      1 självhäftande
      1 självhat
      1 självhjälpsgrupper
      1 självhjälpslitteratur
      1 självhjälpsmetod
      1 självhjälpsmetoder
      1 självhushåll
      3 självhypnos
      1 självidentifierade
      1 självinfektion
      4 självinsikt
      1 själviska
      7 självkänsla
      1 självklar
      1 självklara
      1 självklarhet
      7 självklart
      2 självkontroll
      1 självkontrollen
      1 självkopiera
      2 självläka
      2 självläkande
      2 självläkning
      1 självlärande
      2 självlysande
      1 självmant
      2 självmedicinera
      2 självmedicinerande
      1 självmedicinering
      2 självmedicineringsteorin
      1 självmedvetande
      1 självmedvetandet
      1 självmedvetenhet
      1 självmedvetna
    109 självmord
      1 självmördade
      1 självmördare
      1 självmördaren
      2 självmördarna
      7 självmorden
      1 självmordens
      9 självmordet
      1 självmordhot
      1 självmordnivå
      3 självmordsattack
      2 självmordsattacker
      5 självmordsbenägen
      1 självmordsbenägenhet
      5 självmordsbenägna
      1 självmordsbeteenden
      1 självmordsbombarna
      2 självmordsbrev
      1 självmordsbrigader
     19 självmordsförsök
      4 självmordsfrekvens
      2 självmordsfrekvensen
      8 självmordskris
      1 självmordskriser
      3 självmordsnivå
      1 självmordsnivåerna
      2 självmordsnivån
      2 självmordspakter
      1 självmordsprevention
      1 självmordspreventionen
      2 självmordsrisk
      2 självmordsrisken
      1 självmordssmitta
      1 självmordsstatistik
      1 självmordstal
      5 självmordstankar
      1 självmordstendenser
      1 självmordsuppfattningar
      1 självmordsvåg
      1 självmumifierat
      1 självningssvårigheter
      1 självpåtagna
      1 självpollinering
      1 självrapporterade
      1 självrapportering
      1 självregistrering
      2 självreglerande
      1 självreglering
      1 självrisk
      1 självrisken
      1 självriskerna
      1 självsäkra
      3 självsår
      1 självskada
      5 självskadande
      1 självskadandet
     19 självskadebeteende
      3 självskadebeteenden
      1 självskadebeteendet
      2 självskador
      1 självskattning
      1 självslocknande
      2 självständig
      2 självständiga
      2 självständighet
      8 självständigt
      1 självstimulerar
      1 självstödet
      2 självsuggestion
     16 självt
      1 självtester
      1 självtorka
      6 självuppfattning
      1 självuppskattning
      1 självuppskattningar
      1 självupptagenhet
      4 självvald
      2 självvalda
      1 självvalt
      1 sjärn
      7 sjätte
      5 sjö
     10 sjöar
      1 sjöben
      1 sjöborrar
      1 sjöfarande
      1 sjögräs
      4 sjögrens
      1 sjögurkor
      1 sjöjungfrusyndromet
      1 sjökablar
      1 sjökalkning
      1 sjölök
      1 sjöman
      9 sjömän
      1 sjömännen
      1 sjömärke
      2 sjön
      4 sjönk
      1 sjöräddning
      2 sjörövare
      2 sjösjuka
      1 sjöss
      1 sjövatten
      2 sjöväxter
      1 sjöväxternas
     46 sju
      1 sjua
      1 sjuårsåldern
      1 sjudagars
      1 sjudomar
     37 sjuk
     92 sjuka
     12 sjukan
      1 sjukaste
      1 sjukbesök
    599 sjukdom
    587 sjukdomar
     26 sjukdomarna
      3 sjukdomarnas
      5 sjukdomars
      1 sjukdomde
    659 sjukdomen
     34 sjukdomens
      1 sjukdomepidermoida
      2 sjukdoms
     10 sjukdomsalstrande
      2 sjukdomsalstrare
      1 sjukdomsämnen
      3 sjukdomsbegrepp
      1 sjukdomsbegreppen
      2 sjukdomsbegreppet
      2 sjukdomsbehandlingen
      1 sjukdomsbekämpning
      1 sjukdomsberättelse
      7 sjukdomsbild
     15 sjukdomsbilden
      1 sjukdomsbilder
      1 sjukdomsbilderna
      1 sjukdomsbörda
      2 sjukdomsbördan
      1 sjukdomsdebuten
      3 sjukdomsdiagnos
      1 sjukdomsepisoder
     16 sjukdomsfall
      1 sjukdomsföreteelse
     17 sjukdomsförlopp
     18 sjukdomsförloppet
      1 sjukdomsförlopps
      1 sjukdomsformen
      1 sjukdomsfrågeställningar
      1 sjukdomsframkallade
     11 sjukdomsframkallande
      2 sjukdomsgrupp
      1 sjukdomshistoria
      6 sjukdomsinsikt
      1 sjukdomsinsikten
     10 sjukdomskänsla
      1 sjukdomskategorier
      1 sjukdomsklassifikation
      1 sjukdomslära
      1 sjukdomsliknande
      5 sjukdomsmekanism
      1 sjukdomsmekanismen
      2 sjukdomsmekanismer
      1 sjukdomsmekanismerna
      1 sjukdomsmisstanke
      1 sjukdomsmodellen
      1 sjukdomsmönstret
      1 sjukdomsnivån
      3 sjukdomsorsak
      1 sjukdomsorsaken
      1 sjukdomsorsaker
      2 sjukdomsparanoia
      1 sjukdomsperspektivet
      1 sjukdomsprocess
      2 sjukdomsprocessen
      2 sjukdomsprocesser
      1 sjukdomsprognosen
      1 sjukdomsrelaterad
      1 sjukdomsstadie
      1 sjukdomsstadier
      2 sjukdomsstånd
      1 sjukdomsstarten
      1 sjukdomsstatus
      7 sjukdomssymptom
      1 sjukdomssymptomen
      3 sjukdomssymtom
      1 sjukdomssymtomen
      1 sjukdomssyndrom
      5 sjukdomstecken
      1 sjukdomstecknen
      1 sjukdomstendens
      1 sjukdomstid
      4 sjukdomstiden
     58 sjukdomstillstånd
      5 sjukdomstillståndet
      1 sjukdomstypen
      1 sjukdomsutbrott
      1 sjukdomsutbrottet
      3 sjukdomsutveckling
      7 sjukdomsutvecklingen
      2 sjukdomsyttringar
     34 sjuke
      3 sjukes
      5 sjukförsäkring
      3 sjukförsäkringen
      1 sjukförsäkringsavgift
      2 sjukfrånvaro
      1 sjukfrånvarokostnader
      9 sjukgymnast
      1 sjukgymnasten
      5 sjukgymnaster
      1 sjukgymnastförbundet
     11 sjukgymnastik
      1 sjukgymnastiken
      1 sjukgymnastiska
      1 sjukgymnastutbildningar
      1 sjukhem
      5 sjukhistoria
      1 sjukhistorien
    145 sjukhus
      1 sjukhusapotek
      1 sjukhusbibliotek
      1 sjukhuschefen
      7 sjukhusen
      1 sjukhusens
     24 sjukhuset
      3 sjukhusets
      3 sjukhusfartyg
      3 sjukhusförvärvad
      2 sjukhusförvärvade
      1 sjukhusfysiker
      1 sjukhusfysikerprogrammet
      2 sjukhusinlagda
      3 sjukhusinläggning
      3 sjukhusinläggningar
      1 sjukhusinläggningmedan
      1 sjukhusinskrivningen
      1 sjukhusklinikerna
      1 sjukhusmiljöer
      1 sjukhusmottagning
      1 sjukhusmottagningar
      1 sjukhusområde
      1 sjukhussjuka
      3 sjukhustandläkare
      1 sjukhustandläkarnas
     12 sjukhusvård
      1 sjukhusvården
      3 sjukhusvistelse
      1 sjukhusvistelser
      1 sjukhusyrken
      1 sjukintyg
     16 sjuklig
     11 sjukliga
      1 sjuklighet
      1 sjukligheten
     12 sjukligt
      1 sjukodmen
      1 sjukpenningdagar
      2 sjukplatser
      2 sjukroll
      2 sjukrollen
      1 sjukrollsinnehav
     26 sjuksköterska
      4 sjuksköterskan
      4 sjuksköterskans
      1 sjuksköterskestudenter
      1 sjuksköterskeutbildning
     18 sjuksköterskor
      2 sjuksköterskorna
      1 sjukskriven
      2 sjukskrivningar
      2 sjukskrivningen
      1 sjukstugor
      1 sjukstugorna
      8 sjukt
      1 sjuktransport
     58 sjukvård
      1 sjukvårdande
      5 sjukvårdare
     80 sjukvården
      1 sjukvårdenmedicinen
     11 sjukvårdens
      1 sjukvårdpersonal
      1 sjukvårdsanläggning
      1 sjukvårdsanställda
      1 sjukvårdsartikel
      1 sjukvårdsassocierad
      1 sjukvårdsavgiften
      1 sjukvårdsbefäl
      1 sjukvårdsbehovet
      1 sjukvårdsföretag
      2 sjukvårdsförsäkring
      1 sjukvårdsgrupp
      1 sjukvårdsinrättning
      1 sjukvårdsinrättningar
      2 sjukvårdsinsatser
      4 sjukvårdslagen
      1 sjukvårdslära
      2 sjukvårdsman
      1 sjukvårdsområde
     19 sjukvårdspersonal
      6 sjukvårdspersonalen
      1 sjukvårdsrådgivningen
      1 sjukvårdsspecialist
      1 sjukvårdsstandard
      3 sjukvårdssystem
      4 sjukvårdssystemet
      1 sjukvårdstillstånd
      1 sjukvårdsuppgifter
      2 sjukvårdsupplysningen
      1 sjukvårdsutbildad
      2 sjukvårdsutbildning
      1 sjulingar
      2 sjunde
      7 sjunga
      1 sjungande
      6 sjunger
      9 sjunka
      6 sjunkande
     59 sjunker
      6 sjunkit
      1 sjuttio
      2 sjuttiotalet
      1 sjuttonde
      1 sjutusen
      1 sjvfs
      1 sjvm
    111 sk
      1 �sk
    727 ska
      1 skabb
      1 skabbdjuret
    183 skada
     21 skadad
     35 skadade
      1 skadadedöda
      2 skadades
     37 skadan
      3 skadande
      1 skådande
      1 skadans
     39 skadar
     38 skadas
      1 skådas
      1 skadasymtom
     12 skadat
     10 skadats
      1 skadebegränsning
      1 skadebild
      1 skadechock
     12 skadedjur
      1 skadedjursbekämpare
      1 skadedjursbekämparen
      1 skadedjursbekämpning
      1 skadefall
      3 skadegörare
      1 skadegörarens
      2 skadegörelse
      1 skadeinsekter
      5 skademinimering
      3 skadeområdet
      1 skådeplats
      1 skadeplatsen
      1 skadereducerande
      2 skadereducering
     26 skadereduktion
      1 skadereduktionsåtgärder
      1 skadereduktionsprinciperna
      1 skadereduktionsrörelsens
      3 skaderisken
      1 skådespel
      5 skådespelare
      3 skådespelaren
      1 skådespelarna
      3 skådespelerskan
      1 skadeståndsskyldig
      1 skadevållande
      1 skadeverkan
      3 skadeverkningar
      1 skadeverkningarna
      1 skadjur
     12 skadlig
     47 skadliga
     36 skadligt
    204 skador
     18 skadorna
     13 skaffa
      5 skaffar
      1 skaffat
     10 skaft
      4 skaftade
      1 skaftat
      1 skaftet
      1 skaftlösa
      1 skagerrak
      5 skägg
      1 skäggig
      1 skäggriska
      1 skäggriskan
      1 skäggstrån
      1 skäggstråna
      1 skäggväxt
      1 skäggväxten
      4 skaka
      1 skakade
      3 skakar
      3 skakas
      1 skakiga
      2 skakningar
      1 skäkta
     10 skal
      7 skål
     72 skäl
     30 skala
     11 skalan
      1 skålar
      1 skalas
      1 skalbaggar
      2 skalden
      9 skaldjur
      2 skålen
      6 skälen
      4 skalet
      5 skälet
      1 skålformade
      1 skälig
      1 skäliga
      1 skäligen
    298 skall
      3 skallar
      2 skallarna
      2 skallbasen
      2 skallbasfraktur
      1 skallben
     12 skallbenet
      1 skallbenets
      2 skalle
      1 skallehuvud
     13 skallen
      3 skallens
      1 skallerorm
      1 skallerormsgift
      1 skallform
      1 skallformen
      1 skallfraktur
      1 skallfrakturer
      2 skallighet
      1 skallmissbildningar
      1 skållning
      1 skallskada
      1 skallskador
      4 skällsord
      1 skalltrauma
      7 skalmar
      1 skalmarna
      1 skalömsning
      3 skalor
      1 skalorna
      3 skalpell
      4 skalpeller
      3 skalpen
      1 skalpkylning
      1 skalprotes
      1 skalskydd
      3 skam
      2 skamkänsla
      1 skamkänslor
      1 skamlöshet
      1 skäms
      1 skämtsam
      1 skämtsamt
      3 skandal
      2 skandalen
     12 skandinavien
      5 skandinaviska
      1 skandinaviske
     12 skåne
      3 skånes
      1 skänka
      4 skänkelblock
      2 skänker
      2 skänklar
      1 skänks
      1 skänkte
      1 skannas
      1 skanning
      1 skanningen
      2 skåp
     93 skapa
      8 skapad
     23 skapade
     15 skapades
      1 skapaforma
      1 skapande
      9 skapandet
     52 skapar
      4 skapare
      1 skaparen
     33 skapas
     14 skapat
      6 skapats
      1 skapelse
      1 skapopbandet
      1 skar
      8 skär
      3 skara
     17 skära
      3 skärande
      3 skäras
      2 skärgård
      1 skärklipper
      2 skärm
      1 skärmade
      1 skärmar
      1 skärmarna
     22 skärmen
      3 skärmens
      2 skärmning
      1 skärning
      1 skärningen
      1 skärningspunkt
      1 skaror
      1 skåror
      1 skäror
     14 skarp
      5 skarpa
      2 skärpa
      1 skärpan
      1 skarpare
      1 skärpning
      1 skarpsynta
     10 skarpt
      1 skärpt
      1 skärpta
      1 skärpte
      2 skärptes
      1 skars
      6 skärs
      5 skärsår
      1 skärskada
      1 skärskador
      1 skärskilt
      1 skarv
      1 skärvapen
      1 skarvar
      3 skatta
      6 skattas
      1 skatte
      1 skatteavdraget
      1 skattefinansierad
      1 skattefinansierade
      1 skattehöjning
      1 skatteincitament
      2 skattelättnader
      2 skattemyndigheten
      1 skattemyndigheter
      3 skatter
      1 skattereformen
      1 skatteverket
      2 skattning
      1 skattningar
      1 skattningen
      1 skattningsformulär
      1 skattningsformulären
      1 skattningsskala
      2 skattningsskalor
      1 skattningssystem
      1 skav
      1 skava
      1 skavande
      1 skavanker
      1 skaver
      6 skavsår
    119 ske
      2 sked
      1 skedar
      1 skedarna
     35 skedde
     33 skede
      6 skeden
      2 skedet
      2 skeenden
      1 skeendena
      2 skeletal
      1 skeletala
     23 skelett
      2 skelettben
      1 skelettbesvär
     11 skelettcancer
      1 skelettcancerform
      1 skelettcancerformer
      1 skelettcancerformerna
      1 skelettdeformationer
      1 skelettdestruktioner
      1 skelettelement
     31 skelettet
      4 skelettets
      1 skelettettumören
      1 skelettförändringar
      1 skelettinfektion
      1 skelettinfektioner
      1 skelettlik
      1 skelettmatastaser
      6 skelettmetastaser
      1 skelettmuskelceller
      3 skelettmuskler
      1 skelettmusklerna
      1 skelettmusklernas
      5 skelettmuskulatur
      5 skelettmuskulaturen
      1 skelettmuskulaturens
      1 skelettresorption
      1 skelettrester
      1 skelettröntgen
      1 skelettsegment
      3 skelettskintigrafi
      2 skelettsmärtor
      4 skelettumörer
      1 skelettutveckligen
      2 skelettutveckling
      1 skelettvärk
      1 skellefte
      4 skellefteå
      1 skellefteås
      3 skelning
      1 skelögdhet
      1 skelört
      1 skelörten
      1 sken
      1 �sken
      2 skena
      5 skenan
      1 skenande
      1 skenbar
      6 skenbenet
      2 skenbenets
      2 skendräktighet
      1 skenet
      3 skengraviditet
      3 skenor
      1 skensamband
      2 skepnad
      1 skepp
      2 skepparen
      1 skeppsbesättningar
      3 skeppsbottenfärg
      2 skeppsbottenfärger
      2 skeppskatt
      1 skeppskatter
      1 skeppsråtta
      1 skepsis
      4 skepticism
      1 skeptikern
      2 skeptisk
      1 skeptiska
    374 sker
     39 skett
     12 skick
      8 skicka
      4 skickade
      4 skickades
      1 skickande
     21 skickar
     27 skickas
      2 skickat
      1 skickelig
      1 skicklig
      2 skickliga
      1 skicklighet
      1 skid
      1 skidade
      2 skidåkare
      1 skidbackar
      1 skidfärder
      2 skidspår
      1 skien
      1 skiffer
      1 skiffle
      1 skiffrar
      4 skift
      2 skifta
      7 skiftande
      7 skiftar
      2 skiftarbete
      3 skiftat
      1 skifterna
      1 skiftningar
      1 skiftregister
     15 skikt
      1 skikten
      3 skiktet
      1 skiktets
      1 skiktmetoder
      3 skiktröntgen
      2 skiktsnitt
      1 skild
     23 skilda
      6 skilde
      4 skildes
      4 skildkönade
      1 skildrade
      6 skildrar
      1 skildras
      2 skildrat
      3 skildrats
      1 skildringarna
     51 skilja
      1 skiljaktiga
      1 skiljaktigheter
     14 skiljas
      2 skiljde
      1 skilje
      1 skiljelinje
      1 skiljelinjer
    154 skiljer
      8 skiljs
      1 skiljt
      1 skill
      1 skilld
      1 skillgate
    176 skillnad
     58 skillnaden
     52 skillnader
      1 skillnaderdendriterna
     10 skillnaderna
      1 skills
      7 skilsmässa
      1 skilsmässor
      3 skilt
      1 skimmer
      3 skin
      1 skingras
      1 skinka
      1 skinkan
      1 skinkor
      7 skinkorna
     14 skinn
      1 skinnbaggarna
      6 skinnet
      1 skinnkläder
      1 skinnskorpor
      1 skinnsvampar
      1 skinpick]
      1 [skinpickcom
      1 skinpickcomstoppickingmyskin
      1 skirat
      1 skisserar
      1 skitig
      5 skiva
      3 skivan
      2 skivans
      1 skivas
      1 skivbolag
      1 skivbolaget
      1 skivepitel
     10 skivepitelcancer
      1 skivepitelcancrar
      1 skivepitelet
      1 skivepitelmetaplasi
      1 skivepitelscancer
      1 skivepiteltyp
      1 skivintäkter
      1 skivlingar
     13 skivor
      3 skivorna
      1 skjortor
      1 skjukdom
     11 skjuta
      1 skjutas
      1 skjutbanor
     12 skjuter
      1 skjutklara
      1 skjutning
      1 skjutövningar
      3 skjuts
      2 skjutsa
      9 skjutvapen
      1 skk
      3 skks
      1 sklerodermi
      6 skleros
      1 skleroserande
      3 sklerotier
      6 sklerotierna
      1 sklerotiernas
      1 sklerotiet
      3 sklerotium
      2 sko
      1 sködkörtelrubbningar
      3 skog
      7 skogar
      1 skogarna
      5 skogen
      2 skogs
      1 skogsängar
      1 skogsbingel
      1 skogsbingeln
      1 skogsbrand
      1 skogsbruket
      1 skogsdöende
      1 skogsharar
      1 skogsindustrin
      1 skogslönn
      1 skogsmård
      2 skogsmark
      1 skogssork
      3 skogssorkar
      1 skogssorkarna
      1 skogssorken
      2 skoinlägg
      1 skol
     19 skola
      1 skolad
      4 skolåldern
      1 skolämnena
     35 skolan
      2 skolans
      1 skolår
      1 skolarbete
      1 skolarbeten
      2 skolastikerna
      1 skolbänken
      4 skolbarn
      1 skolbetyg
      1 skolbildning
      2 skolbildningar
      1 skoldagar
      2 sköldberg
      1 sköldbrosk
      1 sköldbroskkannbroskmuskeln
      1 skoldeltagandet
      6 sköldkörtel
      1 sköldkörtelcancer
      1 sköldkörtelenzym
      2 sköldkörtelfunktion
      1 sköldkörtelfunktionen
      3 sköldkörtelhormon
      2 sköldkörtelhormoner
      4 sköldkörtelhormonerna
      1 sköldkörtelhormonreceptorer
     10 sköldkörtelinflammation
     38 sköldkörteln
      8 sköldkörtelns
      1 sköldkörtelproblem
      3 sköldkörtelsjukdom
      1 sköldkörtelsjukdomar
      1 sköldkörtelstimulerande
      1 sköldkörteltillväxt
      1 sköldkörtelvävnad
      1 sköldlöss
      1 sköldpaddor
      1 sköldpaddsskal
      1 sköldskörteln
      1 skole
      1 skolexemplen
      1 skolexemplet
      1 skolfobi
      1 skolform
      1 skolförmåga
      1 skolgång
      1 skolgymnastik
      1 skolhälsovård
      6 skolhälsovården
     14 skolios
      1 skoliosdrabbad
      2 skoliosen
      1 skolioser
      1 skoliosoperation
      1 skoliosopererade
      1 skölj
     12 skölja
      2 sköljas
      1 sköljde
      1 sköljdes
      3 sköljer
      9 sköljmedel
      5 sköljning
      1 sköljningar
      3 sköljningen
      1 sköljningsduscher
      9 sköljs
      1 sköljvätskan
      1 skolkar
      1 skolklassen
      1 skolklasser
      1 skolkning
      2 skolläkare
      3 skolläkaren
      1 skolmassaker
      1 skolmassakrar
      1 skolmatsprogram
      8 skolmedicinen
      1 skolmedicinsk
      2 skolmiljö
      4 skolmiljön
      2 skolning
     14 skolor
      4 skolorna
      1 skolpersonal
      1 skolsituationen
      2 skolsköterska
      1 skolsköterskan
      1 skoltiden
      1 skolundervisning
      1 skolundervisningen
      1 skolungdom
      1 skoluniform
      6 skolvägran
      4 skolvägrar
      1 skolverket
      1 skolverksamheter
      1 skomakaren
      1 skomakartumme
      1 skon
      1 skona
      1 sköna
      1 skonas
      1 sköndals
      5 skönhet
      1 skönheten
      1 skönhets
      1 skönhetsbehandling
      1 skönhetsbehandlingar
      1 skönhetsideal
      1 skönhetsindustrin
      1 skönhetsingrepp
      1 skönhetsinriktade
      1 skönhetsoperation
      1 skönhetsoperationer
      1 skönhetsprodukter
      1 skoningslöst
      1 skönjas
      1 skönlitterära
      3 skönlitteratur
      1 skönlitteraturen
      1 skonsam
      1 skonsamma
      5 skonsammare
      3 skonsamt
      1 skönt
      1 skop
      2 skopa
      1 skopan
      1 skopéa
      6 skopolamin
      1 skoptofil
      1 skoptofila
      2 skoptofili
     16 skor
      3 skör
      5 sköra
      1 skörare
      9 skörbjugg
      2 skörd
      1 skörda
      1 skördade
      2 skördar
      1 skördas
      1 skördat
      2 skördeförluster
      3 skörden
      1 skorna
      1 skorpa
      1 skorpbildning
      1 skorpiongiftödla
      8 skorpiongiftödlan
      2 skorpiongiftödlans
      3 skorpiongiftödlor
      1 skorpiongiftödlorna
      1 skorpionödlan
      1 skorpionödlor
      2 skorpor
      1 skorporna
      1 skorsstenar
      2 skorsten
      1 skorstenar
      1 skorstövlar
      2 skört
      1 skostorlek
      1 skosulor
      2 sköt
      8 sköta
      3 skötare
      1 skötaren
      2 skötas
     17 sköter
      2 sköterska
      1 sköterskan
      9 sköts
      5 skötsel
      1 skötselanvisningen
      1 skötseln
      8 skott
      2 skött
      1 skötta
      1 skötte
      3 sköttes
      1 skottkedja
      4 skottland
      1 skottskada
      1 skotyp
      4 skov
      3 skövde
      1 skövlar
      1 skövling
      1 skovvis
      1 skparietala
      1 skrå
      8 skräck
      1 skräckfilmer
      1 skräckfyllda
      1 skräckhistorier
      1 skräddarjärn
      1 skräddarsydd
      1 skräddarsydda
      1 skräddarsyr
      1 skräddarsys
      1 skrået
      1 skråets
      1 skragge
      1 skrällande
      2 skrämd
      1 skrämda
      1 skrämde
      1 skråmedlem
      1 skrämma
      3 skrämmande
      2 skrämsel
      1 skrämselreflexen
      3 skrån
      6 skräp
      6 skrapa
      1 skrapande
      1 skrapar
      4 skrapas
      4 skrapning
      1 skrapningar
      1 skrapningborstning
      1 skrapsjuka
      1 skratta
      1 skrattar
      1 skråväsendets
      1 skrek
      1 skrep
      1 skreppe
     30 skrev
      1 skrevor
     12 skrevs
      1 skri
      2 skribenter
      1 skrida
      8 skrift
      1 skriftbild
      1 skriften
      9 skrifter
      3 skrifterna
      3 skriftlig
      3 skriftliga
      3 skriftligt
      1 skriftlösa
      1 skriftserier
      9 skriftspråk
      3 skriftspråket
      1 skriftspråkliga
      1 skriftställarna
      1 skriftsystemet
      3 skrika
      1 skriker
     26 skriva
      2 skrivande
      1 skrivandekonsten
     10 skrivas
      2 skrivelse
      7 skriven
     29 skriver
      5 skrivet
      5 skrivförmåga
      2 skrivförmågan
      1 skrivförmågor
      1 skrivhjälpmedel
      1 skrivinlärning
      7 skrivit
      3 skrivits
      3 skrivkramp
      1 skrivmaskinstiden
      8 skrivna
      1 skrivning
      2 skrivpedagogik
     17 skrivs
      2 skrivsvårighet
      1 skrivsvårighetdyslexi
      4 skrivsvårigheter
      1 skrivtecken
      1 skrivutredning
      1 skrivutredningar
      1 skrivutveckling
      1 skrock
      1 skrönor
      1 skrota
      1 skrotning
      1 skrotum
      1 skrov
      7 skrovet
      3 skrovlig
      1 skrubba
      1 skrubbats
      6 skrubbsår
      1 skruden
     15 skrumplever
      2 skrumpna
      1 skrumpnade
      4 skrumpnar
      1 skrupulös
      1 skruv
      1 skruvades
      1 skruvar
      1 skruvpluggar
      1 skruvpluggmassa
      2 skrymmande
      1 skrymseln
      1 skrynkelfritt
      1 skrynklig
      1 skrynklor
      2 skryptorna
      1 skryta
      2 skugga
      3 skuggan
      1 skuggar
      1 skuggig
      1 skuggiga
      2 skuggrika
      1 skuggväxters
     10 skuld
      1 skuldbördor
      2 skulden
      1 skulder
      1 skulderbladet
      3 skuldkänsla
     10 skuldkänslor
      1 skuldra
      5 skuldror
      1 skuldrornas
      7 skull
    409 skulle
      1 skulptera
      1 skulpturala
      1 skulpturerna
      5 skum
      1 skumbehandling
      1 skumcell
      1 skumceller
      2 skumgummi
      1 skumma
      2 skummar
      1 skummet
      1 skumning
      1 skumningen
      1 skumormen
      2 skura
      1 skuren
      1 skurgummeknän
      2 skurit
      1 skurtrasor
      1 skvalen
      1 skvallrar
      7 skvattram
     69 skydd
     72 skydda
     16 skyddad
     15 skyddade
      1 skyddades
     28 skyddande
      1 skyddandet
     47 skyddar
     15 skyddas
      8 skyddet
      1 skydds
      1 skyddsanordningar
      1 skyddsansvariga
      3 skyddsåtgärder
      1 skyddsbågar
      1 skyddsdräkten
      1 skyddsdräkter
      1 skyddsduk
      2 skyddsfaktor
      2 skyddsfaktorer
      4 skyddsglasögon
      1 skyddsgrad
      1 skyddsgud
      1 skyddshandskar
      1 skyddshelgon
      1 skyddshundtjänster
      1 skyddsklass
      1 skyddsklassen
      1 skyddskommittén
      1 skyddsmasker
      3 skyddsmedel
      1 skyddsmekanismer
      1 skyddsnät
      3 skyddsombud
      1 skyddsombuden
      1 skyddsombudens
      4 skyddsombudet
      1 skyddsombudets
      1 skyddsreflex
      1 skyddsrelation
      3 skyddsrond
      1 skyddsronden
      4 skyddsronder
      1 skyddssymbol
      6 skyddsutrustning
      1 skyddsutrustningen
      2 skyddsvakt
      1 skyddsvakter
      1 skyddsvästar
      3 skyddsympning
      1 skyddsynpunkt
      1 skygg
      1 skygghet
      1 skyla
     16 skyldig
      5 skyldiga
      2 skyldighet
      3 skyldigheter
      1 skylla
      1 skyllde
      1 skyller
     47 skylt
      1 skylta
     19 skyltar
      3 skyltarna
     40 skylten
      1 skyltfönster
      1 skymd
      1 skymfar
      1 skymmer
      1 skymning
      1 skymningen
      1 skyms
      1 skymt
      1 skymtats
      3 skynda
      1 skyndsamt
      1 skyskrapa
      2 skyterna
      1 skytiska
      1 skytte
      1 skyttegravar
      1 skyttegravsfeber
      1 skyttegravsfot
     29 slå
      2 släcker
      1 släcks
      2 släckt
      3 sladd
      1 slade
      3 slående
     83 slag
     19 slaganfall
      3 slaganfallet
      1 slagdrabbade
      2 slagen
      1 slaget
      1 slagets
      1 slagfält
      1 slagfältet
      6 slaggprodukter
      3 slagit
      2 slagits
      3 slagminut
      1 slagna
     81 slags
      1 slagverkfamiljen
      2 slagvolym
      1 slaka
      4 slakt
     12 släkt
      2 slaktade
      1 slaktaren
      2 slaktas
      2 släktband
     36 släkte
     11 släkten
      2 släktena
      1 släkter
      1 slakterinäringen
      1 slakteriverksamhet
      1 släkterna
     65 släktet
      1 släktetparvoviridae
      2 släktets
      6 släkting
      9 släktingar
      2 släktingen
      1 släktnamnen
      5 släktnamnet
      2 släktskap
      1 släktstudier
      1 slalom
      5 slam
      3 slamålder
      1 slamålderformula
      1 slamåldern
      1 slamåldrar
      1 slambehandlingen
      1 slambelastning
      1 slambelastningens
      1 slamhantering
      4 slamhanteringen
      1 slamlagret
      1 slamluftning
      1 slammängd
     14 slammet
      1 slammets
      1 slamsvällning
      1 slamvatten
      1 slamvolymen
     15 slang
      1 släng
      2 slänga
      4 slangar
      3 slängas
      1 slängda
      3 slängde
      1 slängdes
      4 slangen
      1 slängen
      1 slangens
      1 slänger
      2 slängs
      1 slängt
      1 slängts
      3 slanguttryck
      1 slankare
      1 slant
      2 släpar
      4 slapp
      1 slappa
     17 släppa
      4 släppas
     34 släpper
      1 slapphet
      1 släppmedel
      5 slappna
     12 slappnar
      1 slappnas
     12 släpps
      2 slappt
      6 släppt
      2 släppte
      5 släpptes
      2 släppts
     34 slår
      2 slarv
      1 slarvat
      1 slarvfel
      4 slarvigt
     15 slås
      1 slash
      5 slåss
      8 slät
      4 släta
      1 slätas
      1 slätbehandling
      1 slätpolerade
      3 slätröntgen
      1 slätröntgenundersökning
      1 slätströk
      4 slätt
      1 slåtterängar
      3 slåttergubbe
      1 slåttergubbeblommans
      1 slåttergubben
      6 slavar
      1 slaveri
      1 slavpojkar
      4 sle
      8 sleep
      1 sleeve
     38 slem
      1 slembarriären
      3 slembildande
      1 slembildning
      1 slemblod
      1 slemfyllda
     27 slemhinna
      1 slemhinnakan
     27 slemhinnan
      1 slemhinnans
      4 slemhinneförändringar
      1 slemhinneinflammation
      1 slemhinnekontakt
      1 slemhinnekörtlar
      1 slemhinnelagret
      1 slemhinnetäckt
      2 slemhinneveck
      1 slemhinneyta
     52 slemhinnor
     30 slemhinnorna
      2 slemhosta
      1 slemliknande
      4 slemlösande
     11 slemmet
      1 slemmig
      1 slemmiga
      1 slemmigt
      1 slemproducerande
      1 slemproduktion
      1 slemproduktionen
      1 slemsäck
      1 slemutsöndring
      1 slet
      1 slicka
      1 slickande
      1 slickar
      1 slickat
      1 slicklapp
      1 slickning
      7 slida
     41 slidan
     14 slidans
      1 slidcancer
      1 slidgången
      2 slidkatarr
      2 slidkramp
      2 slidöppningen
      2 slidsekret
      1 slidväggarna
      3 slinga
      1 slingan
      1 slingorna
      1 slingrande
      2 slingrar
      1 slingrig
      3 slingriga
      1 slinka
      1 slinta
      1 slipad
      1 slipade
      3 slipar
      1 slipas
      1 slipat
      1 sliper
      3 slipning
      9 slippa
     13 slipper
      1 slips
      1 slipsgalge
      1 slipskivor
      2 slirig
      1 slirigare
      4 slita
      3 slitage
      1 slitaget
      1 slitaslängtyp
      1 sliten
      1 sliter
      1 slitet
      1 slitit
      1 slitits
      1 slitkrafter
      1 slitna
      1 slitningsskador
      3 slits
      1 slitsår
      1 slitskadorna
      1 slitstarka
     11 slog
      1 slogs
      2 slöhet
      2 slöja
      1 slöjd
      1 slopeedge
      1 slöseri
      1 slöt
      1 slöts
      1 slott
      1 slottet
      1 slotts
      3 slovenien
      2 slow
      1 slowwave
      3 slu
      1 sluddrigt
      1 slug
      1 sluggish
      5 slump
      2 slumpartat
      2 slumpen
      4 slumpmässig
      1 slumpmässiga
      5 slumpmässigt
      1 slumpvis
      1 slumpvisa
      1 slungade
      5 slungas
      1 slurry
     50 slut
     35 sluta
      8 slutade
      6 slutändan
      1 slutande
     49 slutar
      1 slutarmuskel
      1 slutarökalinjen
      4 slutas
      7 slutat
      1 slutdestinationen
      9 sluten
      1 slutenbilager
      5 slutenvård
      1 slutenvården
      1 slutenvårdsavdelning
     10 sluter
    124 slutet
      2 slutfas
      1 slutfasen
      5 slutföra
      1 slutföras
      1 slutförs
      1 slutfört
      2 slutförts
      5 slutgiltiga
      2 slutgiltigt
      2 slutit
      1 slutlig
      2 slutliga
     48 slutligen
      1 slutligt
      1 slutmål
      1 slutmålet
      1 slutmuskel
      1 slutmuskeln
      8 slutna
      1 slutning
      2 slutningen
      1 slutningsdefekter
      1 slutningshastigheten
      1 slutningstryck
      1 slutparti
      1 slutprodukt
      2 slutprodukten
      2 slutprodukter
      1 slutprodukterna
      2 slutpunkt
      2 slutrapport
      1 slutrapporten
      1 slutrapportens
      1 slutresultat
      5 sluts
      5 slutsats
     23 slutsatsen
     13 slutsatser
      5 slutskede
      4 slutstadiet
      1 slutstenen
      1 sluttermins
      1 sluttningarna
      1 sm
    275 små
      7 småbarn
      1 småbåtshamnar
      1 småbatterier
      1 småbatteritest
      2 småblad
      1 småbladen
      1 småbladens
      1 småbladig
      2 småblåsor
      3 småcellig
      8 småcelliga
      1 smackningar
      1 smådjur
      1 småfåglar
      1 småfisk
      1 småfläckigt
      4 smågnagare
     37 smak
      1 smaka
      2 smakämne
      1 smakämnen
      1 smakämnena
      1 smakande
      7 smakar
      1 smakat
     12 smaken
      3 smaker
      1 smakfattigt
      1 smakförändringar
      1 smakfulla
      1 smakfullt
      2 smaklökar
      1 smaklökarna
      1 småkörtlar
      1 smaksatt
      2 smaksatta
      1 smaksättning
      1 smaksinne
      1 smaksinnerna
      1 smaksinnets
      1 smakuppfattningen
      1 smakupplevelsen
      7 smal
     10 smala
      2 småland
      1 småländska
      1 smalar
      7 smalare
      1 smalarekortare
      1 smalast
      1 smalbandigt
      1 smalben
      1 small
      1 smällare
      1 smallpox
      3 smalnar
      1 smalnas
     11 smalt
      3 smält
      9 smälta
      1 smältas
      2 smälte
      6 smälter
      5 smältning
      9 smältpunkt
      2 smälts
      1 småmängder
     31 småningom
      1 småord
      1 smaragd
      1 smaragdblomma
      7 smärre
      3 smart
      1 smärt
      1 smarta
    198 smärta
      1 smärtadomningarsvaghet
      1 smärtalidandeaffekt
     79 smärtan
      1 smärtanalys
      5 smärtande
      2 smärtaömhet
      1 smartare
      1 smärtattacker
      1 smärtattackerna
      1 smärtbehandlig
      3 smärtbehandling
      1 smärtbehandlingsmetod
      1 smärtbehandlingsmetoderna
      1 smärtbesvär
      2 smärtförnimmelser
      6 smärtfri
      2 smärtfria
      2 smärtfrihet
      5 smärtfritt
      2 smärtgraden
      1 smärtgräns
      2 smärtgränsen
      1 smärthämmande
      1 smärtimpulser
      2 smärtimpulserna
      1 smärtinpulser
      1 smärtkänsla
      3 smärtkänslig
      5 smärtkänslighet
      1 smärtkänslor
      1 smärtkirurgi
     10 smärtlindrande
      1 smärtlindrare
     32 smärtlindring
      1 smärtlindringen
      1 smärtnivå
      1 smärtområdet
     55 smärtor
      3 smärtorna
      1 smärtplåster
      1 smärtreaktion
      1 smärtreaktioner
      4 smärtreceptorer
      1 smärtreceptorernas
      1 smärtretning
     21 smärtsam
      1 smärtsamhet
     17 smärtsamma
     18 smärtsamt
      1 smärtsignaler
      1 smärtsignalerna
      1 smärtskola
     53 smärtstillande
      1 smärtsyndrom
      1 smärtsystemet
      9 smärttillstånd
      1 smärttillståndet
      1 smärttrappa
      4 smärttröskel
      2 småsår
      1 småskador
      1 småskalig
      1 småväxt
      1 småväxta
      1 småvuxenhet
      1 smbg
      2 sme
      1 smear
      1 smeder
      1 smedjanbrygghuset
      8 smegma
      2 smegman
      1 smeka
      1 smekmånadscystit
      1 smeknamn
      1 smeknamnet
      1 smetas
      1 smf
      1 smi
      3 smidig
      1 smidiga
      4 smidigare
      1 smidighet
      3 smidigt
      1 smil
      1 smileys
     12 smink
      1 sminka
      1 sminkade
      1 sminkas
      2 sminket
      1 sminkningstekniken
      3 sminkprodukter
      1 sminksorter
      6 smith
      1 smithfield
      2 smithpapyrusen
      2 smithsonian
     85 smitta
     40 smittad
     61 smittade
     11 smittades
      2 smittagens
      8 smittämne
     17 smittämnen
      4 smittämnena
      6 smittämnet
     68 smittan
     40 smittar
     41 smittas
      1 smittasmittas
     10 smittat
     24 smittats
      2 smittbärande
      6 smittbärare
      2 smittbäraren
      1 smittdosen
      1 smittdosens
      1 smittfasen
      1 smittfri
      1 smittfrihet
      1 smittfritt
      4 smittkällan
      1 smittkällor
      1 smittkedjan
      1 smittkoppa
     51 smittkoppor
      4 smittkopporna
      2 smittkoppsinfektion
      1 smittkoppsutbrott
      3 smittkoppsvaccin
      1 smittkoppsvaccinationen
      2 smittkoppsviruset
      5 smittoämnen
      2 smittoämnet
      1 smittofarliga
      1 smittoförlopp
      1 smittområdet
      1 smittopunkten
      1 smittor
      3 smittorisk
      3 smittorisken
      1 smittorna
      2 smittosamma
      1 smittosamt
      3 smittospridning
      1 smittotecken
      1 smittotillfälle
     13 smittotillfället
      3 smittovägar
      1 smittöverföraren
      2 smittöverföring
      1 smittöverföringen
      1 smittrisk
      1 smittrisken
     44 smittsam
      1 smittsamhet
      3 smittsamheten
     22 smittsamma
      1 smittsammare
      1 smittsammaste
      9 smittsamt
      1 smittsjukdomar
      6 smittskydd
      1 smittskyddinstitutet
      1 smittskyddsinsitutet
     18 smittskyddsinstitutet
      1 smittskyddsinstitutetref
      1 smittskyddsinstitutets
      1 smittskyddsklassade
     21 smittskyddslagen
      4 smittskyddsläkare
      3 smittskyddsläkaren
      1 smittskyddsläkareveterinärer
      1 smittskyddsläkarföreningen
      1 smittskyddsmyndigheten
      1 smittskyddsorgan
      1 smittskyddspliktig
      1 smittspåring
      2 smittspårning
      1 smittspårningsarbetet
      1 smittspårningsåtgärder
      1 smittspårningspliktig
      3 smittspårningspliktiga
      1 smittspridaren
      1 smittspridarna
     17 smittspridning
      2 smittspridningen
      1 smittväg
      3 smittvägar
      1 smittvägarna
      4 smittvägen
      1 smög
      2 smöjning
      1 smokers
      1 smoking
      4 smör
      1 smörblommeväxter
      1 smörets
      1 smörgås
      1 smörgåsar
      1 smörindustrin
      4 smörja
      1 smörjas
      6 smörjer
      3 smörjmedel
      1 smörjningarna
      1 smörjs
      1 smörkullen
      1 smörträden
      1 smsskrivande
      2 smstumme
      1 smuggla
      2 smugglades
      2 smugglas
      1 smugglingen
      2 smula
      1 smulad
      1 smultrontunga
     12 smuts
      1 smutsas
      1 smutsen
      2 smutsig
      4 smutsiga
      2 smutsigt
      1 smutstvätt
      1 smyckade
      2 smycke
      8 smycken
      2 smyckena
      1 smyckerna
      1 smyckesguld
      5 smycket
     10 smygande
      1 smygfilma
      1 smygtittandet
      1 sn
     69 snabb
     40 snabba
      1 snabbar
     56 snabbare
      3 snabbast
      1 snabbaste
      2 snabbhet
      1 snabbmat
      1 snabbökande
      1 snabbsänka
    174 snabbt
      1 snabbtåg
      1 snabbtest
      4 snabbväxande
      7 snabbverkande
      1 snabel
      2 snabeln
      2 snäcka
      3 snäckfeber
      1 snäckfebern
      1 snäckformad
      2 snäckor
      1 snål
      1 snälla
      1 snålskjuts
      1 snapsglas
      3 snar
      2 snår
     57 snarare
     16 snarast
      1 snarkar
      1 snarkljud
     12 snarkning
      1 snarkningar
      2 snarkningarna
      2 snarkningen
      1 snarkoperation
      2 snarlik
      6 snarlika
      1 snarlikt
     41 snart
      1 snäv
      4 sned
      2 snedhet
      1 snedheten
      1 snedtändning
      2 snedtripp
      1 snedvrids
      1 snefyllase
      1 snegla
      2 snett
      1 snetylnmetyl[dimetylaminoetyl]fenylkarbamat
      2 snickare
      1 snickartumme
      2 snickeri
      1 sniffa
      1 sniffandet
      1 sniffning
      1 snigelfeber
      1 sniglar
      1 snille
     40 snitt
      1 snittar
      2 snittbild
      5 snittbilder
      1 snittblommor
      5 snittet
      1 snittöppningen
      6 snö
      1 snöar
      1 snodd
      1 snödroppe
      1 snof
      1 snöigt
      1 snöklädda
      2 snön
      1 snöpa
      6 snor
      1 snörde
      3 snöre
      2 snören
      1 snöret
      1 snörliknande
      2 snörliv
      2 snörlivet
      1 snörning
      1 snorre
      1 snörskenor
      1 snörskoningar
      1 snört
      1 snöstormar
      1 snott
      4 snow
      1 snp
      1 snpmikromatrisanalys
      1 snpmikromatrisanalyser
      1 snreaktion
      1 snurra
      1 snurrande
      7 snurrar
      1 snurrfåtölj
      1 snus
      1 snusa
      1 snusar
      1 snuset
      2 snusnäsdukarna
      1 snut
      1 snutnoja
      1 snuts
      8 snuva
      1 snuvan
      1 snuvig
      1 snygg
      2 snygga
      1 snyggare
      1 snyggt
      2 snyta
      6 so
      2 soap
      1 sobibór
     16 soc
      1 socbegreppet
    103 social
    141 sociala
      1 socialantropologi
      1 socialarbetare
      1 socialbyråer
      1 socialdarwinismens
      1 socialdemokraterna
      1 socialdepartement
      5 socialdepartementet
      1 socialdriftshypotesen
      1 sociale
      1 socialförfattningar
      1 socialförfattningarna
      1 socialförsäkringar
      1 socialförsäkringsminister
      1 socialgrupp
      1 socialgrupper
      1 socialhögskolor
      1 socialhögskolorna
      1 socialhögskolornas
      1 socialidealismen
      1 socialinstituten
      1 socialisationen
      1 socialiseras
      1 socialist
      1 socialistiska
      1 socialkommunal
      2 socialläkare
      1 socialläkaren
      1 socially
     11 socialmedicin
      2 socialmedicinare
      2 socialmedicinarna
      7 socialmedicinen
      2 socialmedicinens
      1 socialmedicinsk
      3 socialmedicinska
      1 socialmedicinskt
      2 socialminister
      1 socialministerium
      1 socialministern
      1 socialministerns
      1 socialnämnden
      1 socialpedagogiskt
      3 socialpolitik
      1 socialpolitiken
      1 socialpolitisk
      4 socialpolitiska
      1 socialpolitiskt
      1 socialpsykiatrin
      1 socialpsykiatriska
      4 socialpsykologi
      1 socialrätt
      1 socialsekreterare
     64 socialstyrelsen
     20 socialstyrelsens
     66 socialt
      4 socialtjänst
      6 socialtjänsten
      2 socialtjänstens
      7 socialtjänstlagen
      1 socialtjänstpolitik
      1 socialutskottet
      1 société
      1 societeten
      1 societetsdamerna
     18 society
      1 socioekomisk
      2 socioekonomisk
      4 socioekonomiska
      1 sociokommunikativt
      2 sociokulturella
      1 sociokulturellt
      2 sociolog
      1 sociologer
     10 sociologi
      1 sociologin
      1 sociologins
      2 sociologiska
      7 socionom
      3 socionomer
      4 socionomexamen
      1 socionoms
      1 socionomutbildning
      2 socionomutbildningen
      1 sociopatbegreppet
      2 sociopati
      1 sockens
      1 sockenstämman
     34 socker
      1 sockeralkoholerna
      2 sockerart
      3 sockerarten
      5 sockerarter
      2 sockerarterna
      1 sockerbitar
      1 sockerbrist
      1 sockerbristen
      1 sockerfri
      1 sockergrupp
      1 sockergruppen
      1 sockerhalt
      1 sockerhalten
      1 sockerhaltig
      1 sockerhaltiga
      2 sockerindustrin
      1 sockerindustrins
      1 sockerintag
      1 sockerkonsumtion
      1 sockerkulör
      3 sockerlag
      1 sockerlagen
      1 sockermängd
      1 sockermolekylerna
      1 sockerrör
      1 sockerrörsodlingar
      1 sockerrörsplantager
      3 sockersjuka
      1 socknar
      1 socknens
      6 sockret
      1 sockrets
      3 soda
      1 sodalösning
     14 söder
      1 söderberg
      1 söderby
      1 söderfalla
      1 söderfaller
      1 södergran
      1 söderhavsljus
      1 söderhavsöar
      2 söderifrån
      1 söderköping
      3 södermanland
      2 södermanlands
      2 södersjukhuset
      1 södertälje
      1 södertörns
      5 söderut
      1 sodoku
      2 sodomi
      1 sodomin
     48 södra
      2 soffa
      1 sofia
      3 sofistikerad
      1 sofistikerade
      1 sofistikerat
      1 soft
      1 sög
      1 sogne
      2 sögs
      2 söhne
      1 soho
      1 soja
      1 sojaallergi
      1 sojabönor
      2 sojamjölk
      2 sojaprodukter
      1 sojaprotein
     50 söka
      7 sökande
      3 sökandet
      3 sökas
      1 sökbar
     60 söker
      1 sökhundar
      1 sökmotor
      2 sökning
      1 soko�owsko
      1 sökorsaken
      3 sokrates
      1 söks
      7 sökt
      3 sökta
      3 sökte
      1 söktjänst
      8 sol
      6 sola
      3 solade
      2 solan
      2 solanaceae
      1 solani
      1 solanin
      4 solanum
      2 solarium
      5 solbad
      1 solbada
      1 solbestrålning
      1 solblekning
      1 solbränd
      1 solbrända
      1 solbrändhetsliknande
      7 solbränna
      1 sold
      4 soldat
     21 soldater
      6 soldaterna
      2 soldaternas
      1 soldaters
     12 solen
      6 solens
      2 solexponering
      1 solfjäder
      1 solfjäderformat
      1 solgel
     13 solglasögon
      1 solglasögonen
      1 solguden
      1 solhatt
      2 solida
      2 solidaritet
      1 solidarpatologien
      1 solider
      1 solig
      2 soliga
      2 soligt
      1 solitärer
      1 solitt
      1 solium
      1 söljor
      1 solkänslig
      4 solkrämer
      1 sollefteå
      1 sollentuna
      1 söllerkollimator
     17 solljus
      1 solljusets
      2 solms
      4 solna
      2 solning
      2 solo
      1 soloinstrument
      1 sololja
      1 sololjor
      1 solosångarens
      1 solrosfrön
      4 solsken
      1 solskydd
      1 solskyddmedel
      1 solskyddsfaktor
      1 solskyddskräm
     11 solskyddsmedel
      1 solskyddsprodukter
      3 solstickan
      1 solstickans
      1 solsting
      1 solstrålar
      1 solstrålarna
      4 solstrålning
      1 solsystemets
      1 soltidabr
      1 solvatisering
  15374 som
      2 soma
      4 somatisering
      1 somatiseringen
      3 somatisk
      7 somatiska
      2 somatiskt
      7 somatoform
      9 somatoforma
      1 somatoformt
      1 somatomediner
      1 somatosensoriska
      5 somatostatin
      1 somatostatinanaloger
      1 somatostatiner
      1 somatostatinet
      1 somatostatinreceptorer
      3 somatotropin
      1 somavert
      1 sombegränsar
      3 someone
      1 somhade
      1 somi
      1 somite
     29 somliga
      3 sömlös
      5 sommar
      2 sömmar
      1 sommaradonis
      1 sommarblomma
      1 sommarblommor
      1 sommardagar
     28 sommaren
      2 sommarfläder
      1 sommargroende
      1 sommarklätt
      2 sommarmånaderna
      1 sömmarna
      1 sommarpälsen
      1 sommarplanteringar
      1 sommarpraktik
      1 sommarvärme
     54 sömn
      7 somna
      1 somnambul
      4 somnambulism
      1 sömnapéer
      1 sömnapne
     26 sömnapné
      6 sömnapnésyndrom
      3 somnar
      1 sömnattack
      4 sömnattacker
      4 sömnattackerna
      3 sömnbehov
      1 sömnbehovet
      5 sömnbesvär
     16 sömnbrist
      2 sömndjup
     32 sömnen
      1 sömnens
      1 sömnepisod
      1 sömnepisodernas
      1 sömnfas
      1 sömnfassyndrom
      1 sömnförlamning
      1 sömnforskning
      2 sömngående
      5 sömngång
      1 sömngångare
      1 sömngångsepisod
      3 sömngivande
      1 sömnhygien
      1 sömnhygienen
      1 sömnhygienråd
      1 sömnig
      1 sömniga
      1 sömnigare
      8 sömnighet
      1 sömnigheten
      1 sömnighettrötthet
      1 sömnklinik
      1 sömnkurer
      1 sömnkvalité
      5 sömnkvalitet
      1 sömnlabb
      1 sömnlaboratorium
      1 sömnlös
     14 sömnlöshet
     10 sömnmedel
      1 sömnmedelsförgiftningar
      1 sömnmedicin
      1 sömnmedicinska
      1 sömnmedlet
      3 sömnmönster
      2 sömnmyokloni
     10 sömnparalys
      2 sömnparalysen
      1 sömnperioden
      1 sömnprat
      8 sömnproblem
      1 sömnrelaterade
      1 sömnrelaterat
      1 sömnrubbningar
      1 sömnrytmen
      3 sömnsjuka
      1 sömnstadier
      1 sömnstadium
      7 sömnstörning
     24 sömnstörningar
      1 sömnstörningen
      1 sömnstudier
      7 sömnsvårigheter
      1 sömntutesläktet
      1 somnus
      1 sömnvanor
      2 somrar
      1 somvisar
     16 son
      1 sonata
      6 sond
      1 sonda
      5 sonden
      1 sonder
     22 sönder
      1 sondera
      1 sönderdela
      3 sönderdelar
      4 sönderdelas
      4 sönderdelning
      2 sönderdelningen
      4 sönderfall
      3 sönderfalla
      2 sönderfallande
      3 sönderfaller
      2 sönderfallskedjor
      2 sönderfallsprodukter
      1 sönderfallsprodukterna
      1 sonderna
      1 sönderskurna
      1 sönderslagna
      1 sondinnehåll
      1 sondmat
      4 sondmatning
      1 sondnäring
      1 sondnäringar
      1 sondnäringen
      1 sondpump
      2 sonen
      7 söner
      2 sonnbyborgström
      1 sönnerdönnes
      3 sonograf
      6 sonografi
      1 sonografiutrustningar
      1 sonographer
      2 sonora
      1 sonoraöknen
      1 sonson
      2 sony
      1 sopa
      1 sopats
      1 sophie
      1 sopis
      1 sopor
      1 soporna
      1 soppa
      1 soppan
      1 soppar
      1 soppo
      1 sopporna
      1 sopransångare
      1 sopranstämma
      1 soprum
      1 soptunnor
      1 soranos
      1 soranus
      2 sorbitol
      1 sorell
     28 sorg
      1 sorgband
      6 sorgen
      2 sorgeprocessen
      5 sorgereaktion
      1 sorgereaktioner
      1 sorgkläder
      2 sorgsen
      1 sorgset
      1 sörja
      4 sörjande
      3 sörjandes
      2 sörjandet
      1 sörjda
      2 sörjde
      3 sörjer
      1 sörjs
      3 sorkar
      1 sorkår
      2 sorkarnas
      1 sorken
      8 sorkfeber
      1 sorkgift
      1 sorkpopulationen
      9 sort
      3 sorten
      7 sortens
     14 sorter
      6 sortera
      3 sorterar
      5 sorteras
      1 sorterat
      1 sortering
      1 sorterna
     51 sorters
      1 sortiment
      3 sortimentet
      1 sorting
     48 sorts
      2 sos
      6 sosfs
      2 sot
      7 söt
      7 söta
      4 sötare
      1 sötat
      1 sötbesk
      1 soten
      1 sotinlagringar
      1 sötma
      3 sötningsmedel
      1 sotos
      1 sötpotatisplantan
      5 sotpunkt
      1 sötsaker
      1 sotspår
      4 sött
      1 sotutveckling
      4 sötvatten
      1 sötvattenskällor
      1 sötvattenssnäckor
      2 sötvattenssniglar
      1 soul
      1 sound
      2 south
      1 southern
      2 soutiengorge
      1 souvenir
      1 souvernirnäsdukar
     21 sova
      2 söva
     12 sovande
      1 sövande
      1 sovandes
      3 sövd
      1 sovdags
     16 sover
      1 söver
      3 sovit
      1 sovjet
      1 sovjeteran
      4 sovjetiska
      6 sovjetunionen
      6 sövning
      1 sövningnarkos
      1 sövningsmedel
      1 sovplats
      1 sovplatser
      1 sovra
      2 sovrum
      1 sövs
      2 sovställning
      5 spa
      1 spaanläggningar
      1 spacer
      1 spaceshipone
      1 späck
      2 späda
      1 spadar
      1 spädare
     37 spädbarn
      3 spädbarnen
      2 spädbarnet
      2 spädbarnets
      3 spädbarns
      1 spädbarnsålder
      1 spädbarnsåldern
      2 spädbarnsdöd
      3 spädbarnsdödlighet
      6 spädbarnsdödligheten
      1 spädbarnsfamiljer
      1 spädbarnsföräldrar
      1 spädbarnshögkonjunktur
      1 spädbarnshuvud
      1 spädbarnskolik
      1 spädbarnsmassage
      1 spädbarnsmassagen
      1 spädbarnsmödrar
      1 spädbarnsmödrars
      1 spädbarnsmord
      1 spädbarnsmortalitet
      1 spädbarnsstadiet
      2 spädbarnstiden
      1 spade
      1 spaden
      2 späder
      1 spadet
      1 spädning
      2 spädningar
      1 spädningsmediet
      1 spädningsproportioner
      2 späds
      1 spain
      1 spainrättning
      2 spaltas
      1 spalter
      1 spalterna
      1 spaltlampa
      2 spaltlampan
      1 spaltningsytor
      1 spån
      7 spänd
      8 spända
      1 spändes
      1 spång
     26 spanien
      2 spaning
      1 spanish
      1 spanjoren
      1 spann
      8 spänna
      1 spännas
      1 spänne
      1 spännen
     12 spänner
      2 spannet
     33 spänning
     19 spänningar
      2 spänningarna
     17 spänningen
      1 spännings
      1 spänningsfältet
      1 spänningsfilm
      1 spänningsförändringar
      1 spänningsförändringen
      4 spänningshuvudvärk
      2 spänningskänsla
      4 spänningskänsliga
      2 spänningsklassningen
      1 spänningsmärkningen
      2 spänningsnivå
      1 spänningsvariationer
     12 spannmål
      2 spannmålen
     10 spannmålsallergi
      1 spannmålsallergier
      1 spannmålspartiklar
      1 spännplatta
      1 spanns
      5 spänns
      1 spännvidd
      1 spansk
     13 spanska
      1 spanskan
      1 spanskspråkiga
      1 spanskt
      1 spänt
      1 spänts
     28 spår
      4 spara
     10 spåra
      1 sparade
      1 sparametrar
      1 sparametrarna
      2 spårämne
      4 spårämnen
      1 sparande
      1 spårande
      1 sparar
      4 sparas
     13 spåras
      1 sparats
      2 spårats
      1 spårelement
      2 spåren
      2 spåret
      1 sparkar
      1 spårmängder
      1 spårområdet
      3 spärr
      5 spärra
      2 spärrar
      1 spärrarna
      1 spärras
      1 spärrblankett
      1 sparrisväxter
      2 sparsam
      5 sparsamt
      1 spartanerna
      2 spårväg
      1 spårvagn
      1 spårvagnar
      1 spårvis
      2 spasm
      6 spasmer
      1 spasmisk
      1 spasmiska
      1 spasmodisk
      1 spasmolytika
      1 spasmolytikum
      1 spasmos
      9 spasticitet
      2 spasticiteten
      7 spastisk
      1 spastiska
      1 spatel
      1 spathulatus
      3 spatial
      3 spatiala
      1 spc
      1 spearman
      1 spearmint
      1 spec
      1 specfika
      3 special
      1 specialartiklar
      1 specialberedda
      1 specialbeställa
      1 specialbeställas
      1 specialdesignad
      4 specialfall
      1 specialfunktioner
      1 specialgud
      1 specialintressen
      1 specialintresserade
      3 specialisera
     11 specialiserad
     22 specialiserade
      2 specialiserar
      3 specialiserat
      6 specialisering
      1 specialiseringsstjänstgöring
      2 specialiseringstjänstgöring
     11 specialist
      1 specialistbehörighet
      1 specialistbeteckningar
      2 specialistbevis
      1 specialisten
      9 specialister
      1 specialisterläkare
      1 specialistexamen
      1 specialistfärdigheter
      1 specialistgren
      1 specialistgrenar
     10 specialistkompetens
      3 specialistläkare
      1 specialistlegitimation
      1 specialistmottagningar
      1 specialistområden
      1 specialistområdet
      1 specialistpsykolog
      5 specialistsjuksköterska
      1 specialisttandläkare
      1 specialisttjänstgöring
      2 specialisttjänstgöringen
      5 specialistutbildad
      3 specialistutbildade
      9 specialistutbildning
      1 specialistutbildningarna
      4 specialistutbildningen
      2 specialistvård
      1 specialistvårdsavdelning
     30 specialitet
      9 specialiteten
      1 specialitetens
     15 specialiteter
      3 specialiteterna
      1 specialitetsindelningen
      1 specialitetsområden
      1 specialkemienheter
      1 specialkliniker
      1 specialkompetens
      1 specialkonstruerad
      1 specialkost
      1 specialkunskaper
      1 specialltillverkas
      1 specialpedagog
      1 specialpedagoger
      5 specialpedagogik
      1 specialpedagogisk
      1 specialpedagogiska
      1 specialregel
      1 specialschampo
      2 specialskolan
      1 specialsolarium
      1 specialstyrkor
      1 specialsydd
      1 specialsytt
      1 specialundervisning
      1 specialutbildade
      1 specialutbildning
      1 specialutformad
      1 specialutformade
      1 specialvarianter
      1 specialversionerna
     44 speciell
     75 speciella
    121 speciellt
      2 species
      1 specificera
      2 specificerad
      3 specificerade
      3 specificerar
      4 specificeras
     10 specificitet
      1 specified
     56 specifik
     87 specifika
      5 specifikation
      2 specifikationer
     57 specifikt
      1 spect
      2 spectrum
      2 speculum
      1 speech
      1 speed
      1 speedad
      1 speedhack
      3 spegel
      4 spegelbild
      3 spegelbilden
      1 spegelbildsvariant
      1 spegelbildsversionerna
      3 spegeln
      1 spegelneuron
      1 spegelneuroner
      3 spegelneuronsystemet
      6 spegelvänd
      3 spegelvända
      2 spegelvändes
      1 spegla
      1 speglande
      4 speglar
      2 speglas
      1 spektra
      2 spektralanalys
      1 spektralfördelning
      1 spektrat
      2 spektrometer
      2 spektroskopiska
     19 spektrum
      4 spektrumanalysator
      4 spektrumanalysatorer
      1 spektrumanalysatorns
      1 spektrumenvelopen
      1 spektrumet
      1 spektrumets
      1 spektrumkomponenter
      1 spekulation
      2 spekulationer
      1 spekulerade
      1 spekulerades
      3 spekuleras
      3 spekulerat
      1 spekulerats
      1 spekulum
     17 spel
     24 spela
      3 spelad
     12 spelade
      1 spelades
      5 spelande
      5 spelandet
     46 spelar
      9 spelare
      1 spelaregrupper
      3 spelaren
      1 spelarens
      1 spelarna
      6 spelas
      5 spelat
      1 spelautomater
      2 spelbanan
     19 spelberoende
      2 spelberoendet
      3 spelen
      4 spelet
      1 spelets
      1 spelfigurer
      1 spelkaraktären
      3 spelmani
      1 spelmiljö
      1 spelmissbruk
      1 spelpjäs
      1 spelplan
      2 spelplanen
      1 spelrelaterade
      1 spelrum
      1 speltvete
      1 spelutvecklare
      1 spelvanor
      1 spematogon
      2 spenar
      1 spencer
      1 spencisternen
      1 spenderade
      3 spenderar
      1 spenderas
      1 spene
      1 spenens
      1 spenkanalen
      1 spenslig
     31 sperma
      2 spermabank
      1 spermabanken
      1 spermabanker
      1 spermadonation
      5 spermadonator
      3 spermadonatorn
      1 spermakvaliten
      3 spermakvalitet
      8 spermakvaliteten
     13 sperman
      1 spermans
      1 spermaproduktionen
      2 spermaprov
      1 spermaticus
      1 spermatogen
      1 spermatogena
      2 spermatogenes
      5 spermatogenesen
      1 spermatogoner
      1 spermatogonier
      1 spermatozioden
      1 spermatozo
      1 spermatozoer
      1 spermavolym
      3 spermicider
     13 spermie
      3 spermieantal
      2 spermieantalet
      1 spermiebildningen
      1 spermiecell
      5 spermiecellen
      3 spermiecellens
      1 spermieceller
      1 spermiedödande
      2 spermiedonation
      1 spermiefunktion
      1 spermiehuvud
      1 spermiekonkurrens
      1 spermiekvaliteten
     19 spermien
      8 spermiens
      2 spermieproduktion
      4 spermieproduktionen
     78 spermier
     41 spermierna
      9 spermiernas
      1 spermiers
      1 spermies
      1 spermietransport
      1 spes
      1 spesialkommando
      1 spetal
      9 spetälska
      1 spetälskan
      1 spetälskekolonier
      9 spets
      1 spetsade
      4 spetsar
      1 spetsbh
     11 spetsen
      1 spetsfot
      2 spetsig
      6 spetsiga
      4 spetsigt
      1 spetskompetens
      1 spetsnazkommando
      1 sph
      2 sphaerotheca
      1 sphenoidale
      1 sphincter
      1 spicata
      2 spice
      1 spieler
      2 spik
      1 spikar
      1 spikböld
      1 spikes
      3 spikklubba
      1 spikklubbor
      5 spill
      1 spilla
      1 spiller
      1 spillet
      3 spillning
      2 spillo
      3 spina
      4 spinal
      1 spinala
      2 spinalanestesi
      6 spinalbedövning
      3 spinalbedövningen
      1 spinalkanalen
      1 spinalnerv
      1 spinalnerver
      1 spinalnerverna
      1 spinalpunktion
      1 spinalvätska
      1 spindelapor
      1 spindelvävsformade
      4 spindelvävshinnan
      1 spindelvävslika
      1 spindelvävslikt
      2 spindlar
      1 spineboard
      3 spineboarden
      1 spineboards
      1 spinigerum
      1 spinn
      1 spinna
      1 spinotalamiska
      1 spiny
      1 spir�a
      5 spiral
      2 spiralct
      6 spiralen
      3 spiraler
      1 spiralfjäder
      1 spiralform
      4 spiralformad
      2 spiralformade
      1 spiralformat
      1 spiralformigt
      5 spiralis
      1 spiralmönstret
      1 spiriller
      1 spirillum
      1 spirit
      1 spiritismen
      1 spirituella
      1 spiroket
      1 spiroketbakterien
      2 spiroketen
      3 spiroketer
      1 spiroketerna
      1 spirometer
      1 spirometrar
      7 spirometri
      2 spirometriundersökning
      1 spironolakton
      2 spirsyra
      1 spis
      4 spisen
      1 spissa
      5 spjälka
      2 spjälkade
      2 spjälkar
     12 spjälkas
      1 spjälkningen
      2 spjälning
      4 spjälor
      2 spjut
      1 spjutformiga
      1 spl
      1 splen
      1 splendens
      4 splenektomi
      3 splenomegali
      1 splints
      1 splitsning
      1 splittras
      1 splittrat
      1 spneumoniae
      1 spokane
      1 spöke
      1 spöken
      7 spola
      1 spolades
      5 spolar
      5 spolas
      1 spole
      1 spolformade
      1 spolierar
      2 spolmask
      1 spolmaskägg
      1 spolmaskangrepp
      1 spolmaskar
      3 spolmasken
      3 spolning
      1 spolvätska
      1 spom
      1 spondartriter
      1 spondylartriter
      6 spondylit
      1 spongiform
      1 spongiforma
      2 sponsorn
      1 sponsrade
      1 sponsras
      1 sponsrat
      2 sponsring
     12 spontan
     13 spontana
      2 spontanabort
      1 spontanaborteras
      3 spontanitet
      1 spontanrapporteringen
     28 spontant
      3 spor
      2 sporadisk
      4 sporadiska
      6 sporadiskt
      1 sporangier
      1 sporangiet
      1 sporangiets
      1 sporangium
      6 sporbildande
      1 sporbildare
      1 sporbildningen
      2 sporen
     25 sporer
      6 sporerna
      1 sporernas
      1 sporform
      2 sporofyten
      1 sporofyter
      1 sporozoiten
      1 sporozoiter
      1 sporozoiterna
      1 sporozoiternas
      1 sporra
      2 sporre
      1 sporren
      1 sporsäckssvampar
      1 sporsäckssvamparna
      1 sporsäcksvamp
      1 sporsäcksvampar
      1 sporsäcksvampen
      1 spörsmål
      9 sport
      2 sportanläggningar
      1 sportar
      1 sportbh
      1 sportdjur
      1 sportdykning
      7 sporter
      1 sportfiske
      1 sporthästar
      1 sportjakt
      1 sportkläder
      1 sportspel
      1 sportutövande
      2 sportutövning
      1 sporulera
      4 spotta
      4 spottar
      1 spottas
      1 spottkobror
      1 spottkörteln
      5 spottkörtlar
      8 spottkörtlarna
      3 spp
     53 språk
      1 språkanvändning
      1 språkbaserat
      6 språkbruk
      1 språkbruket
      1 språkcentrum
      2 språken
     18 språket
      3 språkets
      1 språkfärdigheter
      1 språkförbistringar
      1 språkforskning
      1 språkförståelsen
      2 språkfunktioner
      1 språkfunktionerna
      1 språkhistoria
      1 språkkunskap
     15 språklig
     19 språkliga
      1 språklighet
      2 språkligt
     10 språkljud
      1 språkljuden
      1 språkljudsenheter
      1 språkljudssystemet
      1 språkmönster
      1 språkproduktion
      1 språks
      1 språkstörda
      4 språkstörning
      2 språkstörningar
      1 språkstörningen
      1 språkträning
      5 språkutveckling
      1 språkvårdsnämnd
      1 sprang
      2 språng
      1 sprängämne
      2 sprängämnen
      1 sprängämnesråvara
      1 sprängämnet
      1 sprängas
      1 sprängde
      2 spränger
      1 sprängkraft
      2 sprängmedel
      1 sprängning
      3 sprängört
      1 sprängs
      2 spray
      1 spraya
      1 sprayats
      1 spraybedövas
      1 sprayburk
      1 sprayer
      1 spraying
      1 sprayinhalator
     40 spred
     15 spreds
      3 sprej
      2 spreja
      1 sprejas
      1 sprejburk
      1 sprejen
      1 sprejform
      1 spreta
      1 spretiga
      8 spricka
      1 sprickbildning
     20 spricker
      1 sprickkapslar
      3 sprickor
     61 sprida
      1 spridande
     47 spridas
     19 spridd
     10 spridda
      1 spridde
     55 sprider
     19 spridit
     11 spridits
     84 spridning
     41 spridningen
      1 spridningshistoria
      1 spridningsmetod
      1 spridningsrisk
      1 spridningsrisken
      1 spridningssätt
      1 spridningssättet
      1 spridningsstället
      2 spridningsväg
      1 spridningsvägar
     93 sprids
      6 springa
      1 springande
      7 springer
      4 springmask
      1 springmaskar
      3 springmasken
      3 springor
      8 sprit
      1 sprita
      2 spritdrycken
      3 spritdrycker
      1 spriten
      5 spritt
      3 spritts
      1 spröd
      1 spröda
      1 sprött
      1 sprouting
      1 sprucket
      3 spruckna
      2 sprungna
     13 spruta
      1 sprutade
      2 sprutan
      9 sprutar
     11 sprutas
      1 sprutat
      2 sprutbyten
      1 sprutbytesverksamhet
      1 sprutfobi
      1 sprutkiosker
      1 sprutnålen
     14 sprutor
      2 sprutrum
      1 sprutstick
      2 sprututbyte
      4 sprututbyten
      3 sprututbytesverksamhet
      1 spunnen
      6 sputum
      3 sputumodling
      1 sputumodlingar
      1 sputumprov
      1 spx
      1 spy
      1 spybollar
      1 sq
      1 squash
      2 squeeze
      2 squibb
      4 sr
      1 sramanism
      1 srat
      1 src
      1 srebp
      1 s�rensens
      3 sri
      2 sribosom
      1 srinivasa
      1 srpida
      1 sruta
      2 sry
      1 srygen
      2 srygenen
      1 srys
      3 ss
      1 ßblockerare
      2 ssen
      1 ssf
      2 ssi
      1 ssmän
      2 ssp
      2 sspe
      1 ssr
     11 ssri
      1 ssrier
      1 ssriläkemedel
      1 ssrimedlen
      3 ssripreparat
      1 ssripreparaten
      3 ssrna
      1 �ssrnaviruset
      1 ssrvep
     13 st
      1 sta
     26 stå
     14 stabil
     13 stabila
      2 stabilare
      2 stabilisator
      1 stabilisatorer
      3 stabilisera
      1 stabiliserad
      1 stabiliserade
      1 stabiliserande
      1 stabiliserar
      4 stabiliseras
      2 stabiliserats
      7 stabilisering
      2 stabiliseringen
      1 stabiliseringsbehov
      2 stabiliseringsmedel
      2 stabilitet
      3 stabiliteten
      6 stabilt
      4 stack
      1 stacks
      1 stäcks
     11 stad
      2 städ
      3 städa
      2 städar
      1 städarbetat
      8 städare
      1 städas
      3 städat
     32 staden
      6 stadens
      1 stader
     12 städer
      9 städerna
      2 städernas
      1 städerska
      1 städet
      4 städfirma
      1 städföretag
      2 städföretaget
      4 stadga
      1 stadgades
      1 stadgarna
      4 stadieindelning
     16 stadier
      7 stadierna
     17 stadiet
      4 stadig
      6 stadigt
      1 stadigvarande
     32 stadium
      1 städkvalitet
      1 städmetod
      1 städmetoder
     21 städning
      1 städningen
      2 städpersonal
      2 stads
      1 städsammanhang
      1 stadsdelen
      2 städsegrön
      4 städsegröna
      1 stadsförvaltning
      1 stadshus
      1 stadsjeepar
      1 stadskärnor
      1 stadskarta
      1 stadskrönikören
      1 stadsläkare
      1 stadsmiljö
      1 stadsmiljöer
      1 stadsportarna
      1 stadstrafiken
      1 stadsvakter
      1 städteknik
      1 städutbildningen
     13 stående
      2 staf
      1 stafettläkare
      1 stafylocock
     30 stafylokocker
      3 stafylokockerna
      2 stafylokockinfektioner
      1 stafylokockstam
      1 stag
      1 stagar
      1 stagen
      1 stagnerade
      1 ståhjuling
      1 ståhjulingar
      2 stainback
      1 staket
      1 staketstolpar
     12 stål
      1 stålbladsisättningen
      1 stålcylinder
      1 stålcylindern
      1 stålet
      1 stålets
      1 stålgrå
      1 stålhammar
      1 ståliftar
      1 stalin
      1 stålkonstruktioner
     63 ställa
     23 ställas
      2 ställbar
      4 ställda
      6 ställde
      6 ställdes
     20 ställe
     49 ställen
      1 ställena
     26 ställer
     88 stället
      2 ställföreträdare
     22 ställning
      8 ställningar
      2 ställningen
      2 ställningsfullmakt
      1 ställningsfullmakten
      2 ställningstagande
      4 ställningstaganden
     75 ställs
      2 ställt
      2 ställts
      1 ställverk
      1 stålmannen
      3 stålskenor
      1 stålskodda
      1 stålspets
      1 stålsuturer
      2 stålull
      1 stålyftar
     12 stam
      1 stämband
     26 stämbanden
      5 stämbandens
      2 stämbandscancer
      2 stämbandsförlamning
      2 stämbandsnivå
      2 stämbandspolyp
      1 stämbandsvibration
      2 stämbandsvibrationen
      1 stamberedningen
      6 stamcell
     24 stamceller
      5 stamcellerna
      1 stamcellsbiologi
      1 stamcellsdelning
      1 stamcellsdonation
      1 stamcellsfaktor
      3 stamcellstransplantation
      1 stamcellterapi
      1 stämd
      1 stamhövding
      1 stämläppar
     10 stämläpparna
      5 stämläpparnas
      6 stamma
      4 stämma
      5 stammande
     28 stammar
      3 stammarna
      1 stammat
     12 stammen
      3 stammens
     16 stämmer
     21 stamning
      1 stämningar
      4 stamningen
      1 stamningsbehandlingen
      1 stamningsdagen
      1 stämningsförskjutningar
      3 stämningsläge
      1 stämningslägen
      3 stämningsläget
      1 stämningsstabilisatorer
      1 stamningsterapi
      1 stamningsupplösande
      1 stampfer
      1 stämplade
      1 stämplas
      1 stämpling
      1 stämplingsteori
      4 stämtonslatens
      2 stämtonslatensens
      3 stämvecken
      1 stämveckens
      1 stämvecksförlamning
     13 stånd
      1 ståndaktig
     24 standard
      1 standardavvikelse
      5 standardavvikelser
      1 standardbedövningen
      5 standardbehandling
      1 standardbehandlingen
      1 standarddiagnos
     10 standarden
      3 standarder
      6 standardiserad
     15 standardiserade
      2 standardiserat
      1 standardiserats
      1 standardiserde
      3 standardisering
      1 standardiseringen
      1 standardmetoden
      1 standardmjölk
      1 standardomständigheter
      1 standardpaket
      1 standardpanel
      2 standards
      1 standardsättet
      1 standardsynskärpan
      1 standardterapi
      2 standardtryck
      1 standardvärdena
      1 standardverk
      9 ståndare
      4 ståndarknappar
      1 ståndarknapparna
      7 ståndarna
      1 standartbehandlingen
      1 standartiserade
      2 ståndet
      6 ständig
      4 ständiga
     18 ständigt
      1 ståndort
      1 ståndpunkt
      1 ståndpunkten
      4 ståndpunkter
      1 standvial
      2 stanford
      2 stanfordbinet
      1 stanfordsjukhuset
      1 stanforduniversitetet
      1 stång
      9 stänga
      5 stängas
      3 stängd
      4 stängda
      1 stängde
      2 stängdes
      2 stängel
      2 stängelns
     10 stänger
      1 stänglar
      1 stängningarna
      7 stängs
      1 stängsel
      7 stängt
      1 stängts
      1 stanislav
      2 stank
      1 stänk
      2 stänka
      2 stanken
      1 stanley
     20 stanna
      3 stannade
     23 stannar
      1 stannas
      3 stannat
      1 stansar
      1 stansarna
      1 stapedius
      1 stapediusreflexen
      1 stapes
      1 staphylé
     21 staphylococcus
      1 stapla
      1 staplas
      1 stapylococcus
      2 star
    107 står
     86 stark
     61 starka
     16 stärka
      4 stärkande
     37 starkare
      2 stärkas
      4 starkast
      3 starkaste
      1 starkastora
     15 stärkelse
      1 stärkelserik
      9 stärker
      1 stärkning
      4 stärks
      2 starksprit
    127 starkt
      2 stärkte
      2 stärktes
      1 starlereflexforskningen
      1 starling
      1 starmark
      9 starr
      1 starrbildning
      1 starren
      7 start
     20 starta
     19 startade
     12 startades
     30 startar
      1 startas
      2 startat
      6 starten
      1 startlereflex
      5 startlereflexen
      1 startmolekylerna
      2 startpunkt
      2 startpunkten
      1 startskottet
      1 starttid
      1 stasi
      5 stat
      4 state
     21 staten
     36 statens
     10 stater
      1 staterna
      1 staternas
      1 staters
      5 states
      1 statik
      2 statin
      2 statiner
      1 station
      2 stationär
      2 stationära
      1 stationärt
      1 statisk
      4 statiska
      8 statistical
     33 statistik
      6 statistiken
      1 statistiker
     10 statistisk
     12 statistiska
     16 statistiskt
      6 statlig
     11 statliga
      1 ståtliga
      1 ståtligare
      3 statligt
      4 stats
      1 statsägda
      1 statsbidrag
      1 statsform
      1 statsgemenskap
      2 statskunskap
      1 statsledningen
      1 statslös
      2 statsmedicin
      1 statsmedicinen
      1 statsministern
      1 statssekreterare
      1 statsvetaren
      4 stått
     36 status
      2 statusen
      1 statusmarkering
      1 statusmedvetande
      2 statyer
      8 stav
      4 stavar
      1 stavarna
      2 stavarnas
      5 stavas
      4 stavat
      1 stavelseinitial
      1 stavelsen
      1 stavelser
      1 stavelsermorfem
      1 stavformad
      3 stavformade
      1 stavformat
      1 stavformig
      2 stavformiga
      3 stävja
      1 stavliknande
     15 stavning
      5 stavningen
      1 stavningsprogram
      1 stavningssvårigheter
      1 stavninguttal
      1 steady
      1 stealiten
      1 stearinsyra
      1 steatit
      1 steatos
      1 stefan
     58 steg
      1 stege
      6 stegen
     15 steget
      1 stegförsteg
      1 stegodon
      1 stegomyia
      2 stegrad
      1 stegras
      2 stegrat
      3 stegring
      1 stegringen
      2 stegsvar
      5 stegvis
      1 stein
      4 steiner
      1 steinerhögskolan
      1 steiners
      1 steinkraus
      1 steinman
      1 steins
      1 stekas
      1 stekbord
      1 stekelgift
      3 stekfett
      1 steklar
      5 stekning
      1 stekpanna
      1 stekpincett
      3 steks
      1 stekt
      1 stekyta
      3 stel
      5 stela
      1 stelare
     17 stelhet
      1 stelheten
      1 stelhetstillstånd
      3 stelkramp
      1 stelkrampsbakterien
      1 stelkrampsskydd
      1 stelkrampstoxinet
      1 stellan
      1 stellata
      9 stelnar
      2 stelnat
      1 stelningen
      1 steloperation
      1 stelopererade
      1 stelopereras
      1 stelt
      1 stemcell
     10 sten
     10 stenåldern
      4 stenålderskost
      2 stenålderskosten
      2 stenåldersmänniskor
      1 stenåldersmat
      1 stenansikte
     16 stenar
      1 stenarbetarnas
     14 stenarna
      1 stenarnas
      2 stenbeck
      1 stenbecks
      1 stenbildning
      1 stenbrott
      1 stenbyggandet
      1 stendamm
      2 stendammlunga
      1 stendammslunga
      2 stendhals
      3 stenen
      5 stenenstenarna
      1 stenfrukter
      1 stenfyllning
      1 stenhårda
      1 stenhuggare
      2 steniga
      1 steninsättningar
      6 stenkolstjära
      1 stenkonstruktioner
      1 stenlunga
      1 stenmangeln
      1 stenmurar
      2 stenmurkla
      1 stenolobus
      1 stenophyllus
      6 stenos
      1 stenoser
      1 stenpassion
      1 stenplatta
      1 stenport
      3 stenras
      1 stenristningar
      2 stensalt
      2 stenskott
      9 stent
      1 stenten
      3 stentet
      2 stentoperation
      1 stentyper
      1 stenytan
      1 stephan
      1 stephanie
      2 stephen
      1 stercobilin
      1 stercoralisascaris
      1 stereoisomerer
      1 stereoskopisk
      1 stereoskopiska
      1 stereoskopiskt
      1 stereotyp
      4 stereotypa
      2 stereotyper
      4 stereotypi
     12 stereotypier
      1 stereotypt
      1 stereum
      8 steril
      6 sterila
      1 sterilfas
      4 sterilisera
      3 steriliserade
      4 steriliserades
      4 steriliseras
     17 sterilisering
      2 steriliseringar
      1 steriliseringarna
      1 steriliseringskrav
      1 steriliseringskraven
      2 steriliseringskravet
      1 steriliseringslagsstiftning
      1 steriliseringslagstiftning
     10 sterilitet
      6 sterilt
      1 sterisk
      1 steriskt
      7 stern
      1 sternbergia
      1 sterns
      1 sternum
      1 steroid
      1 steroida
      2 steroidal
      1 steroidbehandling
     22 steroider
      2 steroiderna
      3 steroidhormon
     10 steroidhormoner
      1 steroidhormonproducerande
      1 steroidhormonreceptor
      2 steroidkedjan
      1 steroidprohormon
      1 steroidreceptorer
      1 steroidreglerare
      1 steroidskelett
      1 steroidskelettet
      1 steroidsyntes
     11 stetoskop
      1 stetoskopet
      1 steve
      1 steven
      2 stevenii
      1 stevensons
      1 stewarttreves
      1 steyn
      6 stf
      2 sthöjningsinfarkt
      3 sti
      5 stick
      9 sticka
      2 stickad
     12 stickande
      1 stickas
      1 stickbäcken
      1 sticken
     18 sticker
      3 sticket
      1 stickhål
      1 stickkanalerna
      4 sticklingar
      1 sticklingars
      3 stickmygga
      6 stickmyggan
      3 stickmyggans
      2 stickmyggen
     23 stickmyggor
      5 stickmyggorna
      5 stickmyggornas
      1 stickmyrtenväxt
      1 stickmyrtenväxterna
      4 stickningar
      1 stickningarpirrningarsockerdrickskänsla
      1 stickor
      2 stickprov
      4 sticks
      4 sticksår
      1 sticksåren
      1 stickställe
      1 stickstället
      1 stickvapen
      1 stickverktyg
      2 sticticus
      1 stier
      7 stift
      2 stiftade
      2 stiftelse
      2 stiftelsen
      1 stiftelsens
      3 stiftelser
      1 stiftelserna
      1 stiften
      2 stiftet
      2 stig
     11 stiga
     17 stigande
      2 stigbygeln
     32 stiger
      1 stigit
      1 stigkanter
      2 stigma
      1 stigmatiserad
      3 stigmatiserande
      1 stigmatiseras
      1 stigmatiserat
      1 stigmatiserats
      4 stigmatisering
      2 stigtiden
      4 stil
      2 stilar
      1 stilarna
      1 stilben
      2 stilen
      2 stilförändringar
      1 still
     16 stilla
      2 stillahavsregionen
      8 stillasittande
      6 stillastående
      1 stillbilder
      1 stilleben
      1 stillhet
      1 stillstående
      1 stilnoct
      1 stilnox
      1 stimluans
      1 stimming
     10 stimulans
      1 stimulansen
      1 stimulant
      2 stimulantia
      4 stimulation
      1 stimulationdbs
      2 stimulator
     21 stimulera
      2 stimulerad
      4 stimulerade
      6 stimulerande
     50 stimulerar
     22 stimuleras
      1 stimulerats
     18 stimulering
      4 stimuleringen
      1 stimuleringselektrod
      1 stimuleringssignal
     63 stimuli
     10 stimulit
      8 stimulus
      1 stimulusbegreppet
      1 stimulusen
      1 stimuluset
      1 stina
      2 sting
      1 stinga
      2 stinget
      1 stioxyl
      3 stipler
      2 stiplerna
      3 stirra
      1 stirrar
      1 stituationer
      1 stiumlerar
      2 stjäl
      6 stjäla
      4 stjälk
      9 stjälkar
      3 stjälkarna
      1 stjälkblad
     13 stjälken
      1 stjälkens
      1 stjälpa
      1 stjälps
      1 stjälpt
      1 stjärna
      6 stjärnanis
      1 stjärnanisens
      1 stjärnanisväxter
      1 stjärnformad
      1 stjärnformade
      1 stjärnlikt
      1 stjärnor
      1 stjärnorna
      3 stjärten
      1 stk
      1 stläkare
      1 stläkaren
      1 stockad
      1 stockade
      1 stockar
     55 stockholm
      1 stockholmföretaget
     22 stockholms
      1 stockholmsbaserade
      1 stockholmsområdet
      1 stockholmsreglementet
      2 stockholmssyndromet
      4 stockholmstrakten
      1 stockholmsutställningen
      3 stockningen
     26 stod
    116 stöd
      1 stödbehandling
      1 stödblad
      1 stödd
      1 stödde
      2 stöddes
      7 stöder
      6 stödet
      3 stödfunktioner
      1 stödgrupper
      1 stödinsatser
      8 stödja
      9 stödjande
      1 stödjeceller
      1 stödjemedel
     10 stödjer
      2 stödjevävnad
      1 stödjevävnader
      1 stödjs
      1 stödpunkter
      1 stödrör
      6 stöds
      1 stödskenan
      1 stödskenor
      1 stödstrumpa
      2 stödstrumpor
      1 stoet
      1 stoffurval
      1 stoft
      2 stokastisk
      1 stökigt
      1 stökiometrisk
      3 stol
      2 stolar
      2 stolarna
      3 stöld
      3 stölden
      1 stölderna
      1 stöldgodset
      1 stöldskydd
      1 stöldskyddsföreningens
      4 stolen
      2 stolgången
      1 stolpar
      5 stolpiller
      2 stolpillret
      1 stolsrygg
      2 stolt
      1 stolta
      1 stolthet
      1 stoltsera
      2 stoma
      1 stomatis
      1 stomatit
      1 stomatologi
     12 stomi
      1 stomibandagestomipåse
      1 stomibandaget
      7 stomin
      1 stomins
      3 stomioperation
      1 stomioperationen
      1 stomipatient
      1 stommen
      1 ston
      1 stone
      3 stop
      2 stopette
      1 stopkonfekt
     14 stopp
     25 stoppa
      1 stoppad
      1 stoppades
      8 stoppar
     12 stoppas
      1 stoppat
      3 stoppet
      1 stopplatta
      2 stopplikt
      1 stoppning
      1 stoppningsrätt
      1 stöpt
    445 stor
     20 stör
    443 stora
      7 störa
     12 störande
      5 störas
     82 storbritannien
      2 storbritanniens
      1 storbröstade
      2 storbystade
     37 störd
      5 störda
      1 störde
      1 stördes
      5 store
      1 störfiskar
      1 storformat
      1 storformatskameror
      2 storfothöns
      1 storhet
      1 storheten
      3 storheter
      2 storheterna
      1 storhetstid
      4 storhetsvansinne
      3 storhjärna
      8 storhjärnan
      1 storhjärnsanlagets
      1 storhushåll
      1 storkok
      1 storkök
     99 storlek
     18 storlekar
      1 storlekarna
     26 storleken
      2 storleksacceptans
      1 storleksförändring
      1 storleksklassen
      1 storlekskontroll
      1 storleksökningen
      1 storleksordning
      8 storleksordningen
      1 storleksskillnad
      1 stormades
      1 stormaktstiden
      2 stormarknaderna
      3 stormavdelningarna
      1 stormhatt
      2 stormhattssläktet
      1 stormning
      1 stormördare
    120 störning
    171 störningar
     14 störningarna
      1 störningarnas
      1 störningars
      1 störningarsjukdomstillstånd
     32 störningen
      1 störra
    408 större
      1 störreodlade
     12 störs
      1 storsäljare
      1 storskalig
      2 storskaliga
      1 storskaligt
     44 störst
    172 största
      1 storstaden
      1 storstäder
      2 storstäderna
      4 storstädning
      1 storstadsfenomen
      1 storstadsområdet
      1 störste
    205 stort
      1 stört
      1 störta
      2 stortå
      1 störtades
      1 stortampn
      8 stortån
      1 storväxt
      1 storväxta
      1 storvuxna
      1 story
      3 stöt
      5 stöta
      1 stötande
      6 stötar
      3 stötas
      1 stötdämpande
     12 stöter
      1 stötkänsligt
     12 stöts
      1 stötta
      1 stöttade
      1 stöttande
      1 stöttepelare
      1 stötvågsbehandling
      1 stötvågslitotripsi
      4 stövsländor
      1 stövsländorna
      1 strabon
      5 sträck
      8 sträcka
      2 sträckan
      1 sträckbänk
     26 sträcker
      1 sträckmetall
      1 sträckmetallcylinder
      3 sträckning
      2 sträckningen
      6 sträckor
      4 sträckreceptorer
      1 sträckreflex
      2 sträckreflexen
      3 sträcks
      4 sträckte
      1 straet
     18 straff
      1 straffad
      4 straffades
      1 straffansvar
      1 straffar
      2 straffarbete
      2 straffas
      2 straffbart
      1 straffbelagt
      5 straffet
      1 straffkompanier
      2 strafflagarna
      1 strafflagstiftningen
      2 strafflöst
      1 straffmyndig
      1 straffrättsligt
      1 straffspark
      1 straffvärde
      1 straffyrkandet
      2 strahlenschutz
      1 straits
      1 stråk
      1 stråke
      1 strål
      3 stråla
      1 strålande
     13 strålar
      1 strålarnas
      1 strålbärarna
      2 strålbehandlas
      1 strålbehandlig
     43 strålbehandling
      1 strålbehandlingar
      3 strålbehandlingen
      1 strålbehandlingsavdelningarna
      2 strålbehandlingsavdelningen
      1 strålbehandlingsmaskin
      1 strålbehandlingspersonalen
      1 strålbehandlingsplanen
      1 strålbehanlding
      1 strålblommor
      2 stråldesinfektion
     10 stråldos
      9 stråldosen
      3 stråldosens
      8 stråldoser
      1 stråldoserna
      4 stråle
     10 strålen
      2 strålens
      1 strålfält
      1 strålfältet
      1 strålforskning
      1 �strålframdrivning
      1 strålfysikalisk
      1 strålgången
      6 strålkälla
      5 strålkällan
      1 strålkällankällorna
      9 strålkällor
     22 strålkällorna
      3 strålkällornas
      1 strålkänsligheten
      1 strålkastarbelysning
      1 strålkirurgi
      1 strålknippe
      1 strålkroppen
     93 strålning
      1 �strålning
      2 strålningar
     30 strålningen
      1 strålningens
      1 strålningsbehandling
      3 strålningsbiologi
      2 strålningsenergi
      1 strålningsexponering
      1 strålningsflöde
      1 strålningsfri
      1 strålningsfria
      7 strålningsfysik
      1 strålningsgraden
      1 strålningsnivå
      1 strålningsnivåer
      1 strålningsonkologer
      1 strålningsrisk
      1 strålningsriskerna
      1 strålningssjuka
      1 strålningsskador
      1 strålningsterapeutisk
      2 strålningstyp
      1 strålningstypernas
      1 strålningsutrustning
      2 strålreaktioner
      1 strålsäkerhet
      1 strålsäkerhetsmyndigheten
      1 strålsäkerhetsmyndighetens
      2 strålsjuka
      3 strålskydd
      1 strålskyddsarbetet
      1 strålskyddsinstitut
      2 strålskyddssammanhang
      1 strålslag
      1 strålspärr
      1 strålterapi
      1 strålterapin
      4 strama
      2 stramar
      1 stramas
      3 stramonium
      1 strån
      7 strand
      1 strandade
      2 stranden
      5 stränder
      2 stränderna
      1 strandhäll
      1 strandkanten
      1 strandkanter
      1 strandkärr
      7 strandvial
      4 sträng
      4 stränga
      3 strängar
      1 strängare
      1 strängarna
      1 strängarnas
      1 strange
      3 strängen
      2 stränginstrument
      1 strängnäs
      4 strängt
      5 strasbourg
      1 strassburg
      1 strategi
     20 strategier
      1 strategin
      1 strategisk
      3 strategiska
      1 stratosfären
      2 stratum
      2 strauss
      1 straussglass
      2 sträv
      3 sträva
      8 strävan
      6 strävar
      1 strävhårig
      1 strävhåriga
      2 strävhet
     36 strax
      1 streching
      9 streck
      1 strecken
      1 strecket
      1 streckgubbe
      1 stred
      4 street
      1 strep
      1 strepsils
      1 streptavidin
      1 streptobacillus
      1 streptococcal
     11 streptococcus
      2 streptokock
      2 streptokockarter
     26 streptokocker
      7 streptokockinfektion
      1 streptokockinfektionen
      4 streptokockinfektioner
      3 streptomyces
     28 streptomycin
    182 stress
      2 stressa
      3 stressad
      3 stressade
      4 stressande
      1 stressaxel
     15 stressaxeln
      3 stressaxelns
      1 stressbehandling
      1 stressbelastning
      1 stressboll
      7 stressen
      1 stressfaktor
      1 stressfaktorer
      2 stressfraktur
      3 stressfrakturer
      1 stressfull
      1 stressfylld
      1 stressfyllda
      1 stresshantering
      1 stresshormon
      5 stresshormoner
      2 stresshormonerna
      2 stresshormonet
      1 stressjukdom
      1 stresskänslor
      1 stresslösande
      1 stressmage
      1 stressmoment
      1 stressmuskeln
      6 stressor
      1 stressoren
     24 stressorer
      7 stressorerna
      8 stressreaktion
      3 stressreaktioner
      1 stressreaktionerna
      4 stressreduktion
      1 stressreglering
      1 stressrelaterad
     10 stressrelaterade
      1 stressrelaterat
      1 stressresponser
      1 stress�sårbarhetsmodellen
      1 stresstillstånd
      1 stressutlöst
      1 stressutlösta
     13 stressyndrom
      1 stressystem
      1 stretcha
      3 stretching
      1 stretchningsövningar
      1 stretchreceptorer
      7 striae
      1 striatal
      2 striatum
     12 strid
      3 strida
      4 stridande
      2 striden
      2 strider
      2 striderna
      1 stridor
      1 stridsfordon
      1 stridsgrupper
      5 stridsmedel
      1 stridspiloter
      1 stridssjukvårdare
      1 stridsskrift
      1 stridssystem
      1 stridströtthet
      4 stridsutmattning
      1 stridsutmattningen
      1 stridsvagnars
      1 stridsvagnskanoner
      1 striglas
     22 strikt
     13 strikta
      1 striktare
      1 striktur
      1 strikturbildningar
      1 strikturer
      1 strilande
      1 strimlar
      1 strimlas
      1 strimlorspån
      2 strimmor
      1 stringanpassad
      1 stringenta
      1 stringtrosor
      1 striptease
      1 strix
      1 ströas
      1 strobilation
      4 stroboskop
      2 stroboskopet
      5 strödda
      1 strofantsläktet
     78 stroke
      1 strokedrabbade
      1 strokeenhet
      1 strokeförbundet
      1 strokekampanj
      1 stroken
      1 strokepatienter
      1 strokerehabilitering
      1 strokesjukvård
      2 stroketeam
     16 ström
      4 stroma
      1 stromacell
      2 stromaceller
      1 stromacellerna
      1 stromacellstumör
      1 stroman
      1 stromaskikt
      1 stromat
      1 strömbäck
      1 strömbad
      1 strömbrytare
      2 stromeyer
      2 strömförsörjning
      1 strömförstärkningsfaktor
      2 strömma
     20 strömmar
      1 strömmatning
      8 strömmen
      2 strömning
      2 strömningen
      1 strömstöt
      2 strömstyrka
      2 strömstyrkan
      2 strongyloides
      3 strontium
      1 strontiumklorid
      1 strophanthus
      1 strophion
      1 strophium
      1 strös
      1 strösocker
      1 strövstigar
     65 struktur
      1 strukturalistisk
      1 strukturändring
      1 strukturbestämdes
      1 strukturdynamik
      2 strukturell
      4 strukturella
      6 strukturellt
     18 strukturen
      1 strukturens
     37 strukturer
      2 strukturera
      2 strukturerad
      3 strukturerade
      1 strukturerar
      2 struktureras
      3 strukturerat
      5 strukturerna
      1 strukturförändring
      1 strukturförändringar
      1 strukturförändringen
      1 strukturformeln
      1 strular
     10 struma
      2 strumpa
      3 strumpor
      1 strumporna
      3 strunta
      2 struntar
      1 strupe
      6 strupen
      2 strupens
      3 struphuvud
     23 struphuvudet
      4 struphuvudets
      3 struplocket
      1 struplockets
      1 strupreflexen
      1 strutade
      1 strychnos
      1 stryk
      2 strykas
      3 stryker
      9 strykjärn
      2 strykjärnen
      2 strykjärnet
      2 strykjärnets
      3 stryknin
      2 strykning
      1 strykningar
      1 strykpressa
      2 stryks
      1 stryktålig
      1 stryparsjukan
      2 stryper
      3 stryps
      2 ststräcka
      1 ststräckan
      4 sttjänst
      2 stubbar
      1 stubbdyna
      1 stubbdynan
      1 stubbdynsvampen
      1 stubben
      1 stubin
      3 stucken
      1 student
      6 studenter
      1 studenterna
      2 studentlägenheter
      2 studentlitteratur
      1 students
     46 studera
      1 studerad
     17 studerade
      3 studerades
      1 studerande
     24 studerar
      1 studerarbr
     29 studeras
     16 studerat
      8 studerats
    131 studie
      1 studieår
      1 studiedeltagare
      1 studieframgångar
      2 studiegång
      1 studiegången
      1 studiegrupperna
      1 studiemedel
     39 studien
      3 studiens
      2 studieobjekt
      1 studieplatser
      1 studieprotokoll
    281 studier
     13 studierna
      1 studiernas
      2 studiers
      1 studier[vilka]
      5 studies
     15 studiet
      2 studieteknik
      1 studietekniken
      1 studietiden
      1 studioalbum
      1 studiobelysningen
      1 studion
      1 studior
      1 studium
      1 studsande
      1 studsar
      5 study
      1 stuff
      1 stuga
      1 stuider
      2 stukning
      1 stum
      1 stumfilmseran
      1 stumfilmsstjärnor
      2 stumhet
      1 stumma
      1 stumpen
      2 stumt
     12 stund
      3 stunden
      1 stundens
      2 stunder
      3 stundom
      1 stunds
      2 stundtals
      1 stungen
      1 stungna
     14 stupor
      2 stuporn
      1 stupur
      2 sturgewebers
      1 sturlason
      2 stussen
      1 stuttgart
      1 styckat
     12 stycke
     27 stycken
      2 stycket
      2 styckl
      1 styfninsyra
      2 stygn
      1 styloglossus
      1 stympande
      1 stympning
      1 stympningar
      1 styng
      1 styngets
      1 styngfluga
      3 styngflugor
     33 styr
     15 styra
      3 styrande
      2 styras
      2 styrd
      1 styrda
      2 styrdes
      1 styre
      4 styrelse
      4 styrelsen
      1 styrelseordförande
      1 styrelser
      1 styren
      1 styrenplast
      2 styret
      1 styrgrupp
      1 styrhytter
      1 styrjärn
     32 styrka
      5 styrkan
      2 styrke
      1 styrkeprov
      1 styrker
      1 styrketräning
      2 styrkor
      2 styrkorna
      1 styrks
      1 styrkula
      1 styrleder
      1 styrlist
      2 styrning
      1 styrningen
      1 styrplatta
      1 styrpunkt
      1 styrpunkter
     37 styrs
      1 styrspak
      2 styrspakar
      1 styrstång
      2 styrt
      1 styrts
      1 styrutrustningen
      2 styva
      1 styvare
      2 styvhårig
      3 styvhet
      2 styvnar
      1 su
      3 subakut
      2 subakuta
      1 subandinus
      4 subarachnoidalblödning
      5 subaraknoidalrummet
      1 subdermal
      1 subendokardiell
      1 subenheten
      4 subenheter
      1 �subenheter
      4 subenheterna
      1 subenhetsvacciner
      1 subfertilitet
      1 subfornikala
      1 subgingival
      4 subglottala
      4 subglottalt
      2 subject
      1 subjekt
      1 subjekten
      5 subjektet
      7 subjektiv
      5 subjektiva
      3 subjektivt
      1 subklinisk
      2 subkliniska
      1 subkomissurala
      3 subkortikala
      3 subkultur
      1 subkulturer
      8 subkutan
      3 subkutant
      1 sublimerar
      1 sublimeras
      4 sublimering
      2 sublingual
      1 sublinguala
      1 sublingualis
      2 subluxationer
      1 submaximalt
      1 submission
      1 suboptimal
      1 suboptimala
      1 subq
      8 subsahariska
     16 subsp
      1 subspecialiteter
      1 substances
     54 substans
      3 substansberoende
      2 substansdroger
      1 substansdrogshistorik
     61 substansen
      2 substansens
     71 substanser
      5 substanserna
      1 substanservävnader
     10 substansmissbruk
      3 substansrelaterade
      1 substituerad
      9 substitut
      1 substituteras
      1 substitutet
      3 substitution
      1 substitutionsbehandling
      2 substitutionsreaktion
      1 substitutionsreaktioner
      3 substrat
      1 substratet
      3 subtil
      4 subtila
      1 subtilis
      1 subtrahera
      1 subtraheras
      5 subtropiska
      1 subtyp
      5 subtypen
     10 subtyper
      1 subtyperna
      1 subulatus
      2 subutex
      1 subvention
      1 subventionerade
      1 subventionerar
      1 subventionssystemet
      1 subventrikulära
      5 succé
      2 succén
      1 success
      1 succession
      2 successiva
     27 successivt
      2 succinylcoa
      1 succubus
      1 suck
      1 sucking
      4 suckulenta
      1 suda
     11 sudan
      3 sudarium
      1 suddig
      1 suddiga
      2 suddigt
      1 suecica
      1 suffix
      1 sufism
      1 sufismen
      2 sug
     21 suga
      4 sugande
      1 sugas
      2 sugdränage
      1 sugeffekt
     12 suger
      1 suget
      1 sugförmåga
      1 sugga
      1 suggan
      1 suggererats
      4 suggestion
      1 suggestioner
      1 suggestiva
      1 suggor
      4 sugit
      1 sugits
      1 sugklockan
      1 sugkoppor
      4 sugmaskar
      1 sugmasksläktet
      2 sugning
      1 sugningen
      1 sugorgan
      7 sugs
      1 sugskålar
      1 sugsnabel
      1 sugsnabeln
      2 sugtablett
      3 sugtabletter
      1 sugtrådar
      3 suicid
      1 suicida
      1 suicidal
      1 suicidala
      3 suicide
      1 suicidförsök
      1 suicidologi
      1 suicidprevention
      1 suicidrisk
      1 suicidrisken
      1 suisse
      4 sula
      1 sulan
      1 sulcus
      1 sulfa
      1 sulfas
      1 sulfatderivat
      1 sulfatet
      1 sulfatgrupper
      1 sulfatprocessen
      1 sulfidmalm
      1 sulfitprocessen
      2 sulfonamid
      1 sulfonamiden
      1 sulfonamidens
      3 sulfonamider
      1 sulfonamidresistens
      1 sulforafan
      1 sulformig
      1 sullivan
      1 sulorna
      1 sulphureus
      1 sultan
      1 sum
      1 sumac
      1 sumak
      2 sumakväxter
      2 sumer
      1 sumererna
      2 sumeriska
      7 summaformel
      5 summaformeln
      1 summan
      1 summary
      1 summer
      3 summera
      1 summeras
      1 summor
      1 sumpfeber
      1 sumpsnäcka
      2 sun
      1 sunburn
      1 sund
      2 sunda
      2 sunday
      1 sundby
      1 sundell
      1 sundhetskollegium
      1 sundstedt
      2 sundsvall
      1 sungai
      1 sungais
      2 sunlight
      1 sunnaas
      1 sunstar
      3 sunt
      1 suntan
      1 suominen
      6 super
      1 superfertilisation
      1 superheterodyntekniker
      1 supérieure
      1 superinfektion
      7 superior
      1 superiora
      1 superiort
      1 superklar
      1 superkompensera
      1 superkomspensation
      1 superlim
      2 superlimmet
      1 supermodell
      1 supernovor
      1 superoxidradikaler
      1 superstars
      2 supervising
      1 supply
      3 support
      1 supporting
      1 suppositoriet
      1 suppositorium
      1 suppression
      1 suppressiontestet
      1 suppressorgen
      3 suppressorgener
      1 supragingival
      1 supraledande
      1 supramolekylär
      1 supraoptiska
      2 suprapubisk
      1 suprarenales
      1 supraventrikulär
      2 supraventrikulära
      2 sur
     18 sura
      2 surare
      1 surditas
      1 sure
      3 surfaktant
      1 surfning
      2 surgery
      3 surhetsgrad
      1 surhetsreglerande
      1 surmafolket
      1 surra
      1 surrealister
      1 surrogatmamma
      1 surrogatmamman
      1 surrogatmodern
      1 surrogatmödraskap
      6 surt
      1 survivor
      4 susan
      1 susande
      1 susceptibilitet
      2 sushi
      5 sushruta
      2 sushrutas
      1 susningar
      3 suspectum
      6 suspension
      2 suspensioner
      1 susruta
      1 suszo
      1 sutra
      4 sutras
      6 suttit
      4 sutur
      1 suturen
     26 suturer
      4 suturerna
      1 suturknut
      1 suturnålar
      1 suturtillverkare
      1 suturtrådar
      1 suturtråden
      1 suzuki
      6 sv
      1 sva
     29 svag
     14 svaga
     18 svagare
      3 svagbegåvade
      2 svågen
     27 svaghet
      4 svagheter
      1 svaghets
      1 svaghetstillstånd
      1 svågor
      1 svagström
     36 svagt
      1 sval
      5 svala
      1 svalare
      1 svald
      2 svalda
      1 svalde
     18 svalg
     37 svalget
      2 svalgets
      1 svalginfektion
      1 svalgmuskulaturen
      1 svalgprov
      1 svalgregionen
      1 svalgringen
      1 svalgrummet
      1 svalgtonsillen
      1 svälj
     18 svälja
      4 sväljer
      8 sväljning
      7 sväljningen
      2 sväljningsreflexen
      3 sväljningsstörningar
      5 sväljningssvårigheter
      1 sväljningssvårigheterna
      2 sväljprocessen
      1 sväljreflex
      3 sväljs
      3 sväljsvårigheter
      2 svalka
      2 svalkar
      1 svalkas
      9 svälla
      7 sväller
      2 svällkroppar
      7 svällkropparna
      2 svällkroppen
      1 svällkroppsvävnad
      1 svalna
      1 svalört
      7 svalt
     18 svält
      4 svälta
      1 svältande
      1 svälten
      1 svältketoner
      1 svältoffer
      1 svältrelaterade
     38 svamp
      1 svampangrepp
     52 svampar
      3 svamparna
      7 svampart
      2 svamparter
      1 svampböcker
      1 svampboll
      1 svampbollar
      1 svampdjur
      2 svampdödande
     37 svampen
     14 svampens
      1 svampfloran
      4 svampförgiftning
      1 svampgifter
      1 svampgrupper
      1 svampiga
     11 svampinfektion
      5 svampinfektioner
      1 svampkropp
      5 svampmeningit
      1 svamporganismer
      1 svampplockare
      1 svampplockning
      1 svamprelaterad
      1 svampriket
      2 svampsjukdom
      1 svampsjukdomar
      1 svampsporerna
      1 svan
      1 svanborg
      1 svanen
      4 svänga
      1 svängande
      5 svänger
      1 svängning
      8 svängningar
      2 svängningarna
      1 svängningsmaximum
      1 svängt
      1 svank
      2 svankrygg
      9 svans
      2 svansar
     11 svansen
      2 svanskotan
      1 svanstipp
      1 svante
     52 svar
    150 svår
      7 svara
    153 svåra
      5 svarade
      1 svarande
     46 svarar
     67 svårare
      3 svårartad
      2 svårartade
      3 svarat
      1 svårbedömda
      1 svårbegriplig
      1 svårbegripligt
      3 svårbehandlad
      3 svårbehandlade
      1 svårbehandlat
      1 svårbemästrade
      1 svårbestämbar
      5 svärd
      1 svärdbärare
      1 svårdiagnosticerat
      2 svårdiagnostiserad
      1 svärdssmeder
      1 svaren
      6 svaret
      1 svårgripbara
      1 svårhanterat
     21 svårighet
      3 svårigheten
     76 svårigheter
     11 svårigheterna
     12 svårighetsgrad
      3 svårighetsgraden
      5 svårighetsgrader
      1 svårighetsgraderna
      1 svårjoniserat
      1 svårjusterat
      1 svårkontrollerbara
      7 svårläkta
      4 svårlöslig
      2 svårlösliga
      3 svårlösligt
      1 svärmande
      1 svärmiska
      2 svårmod
      1 svårnedbrytbara
      1 svårnedbrytbart
      3 svårodlad
      1 svarsalternativ
      1 svarsandel
      1 svarsfrekvens
      1 svarsfrekvensen
      1 svårsmält
      1 svårstuderad
      1 svårstuderade
     41 svart
    199 svårt
     26 svarta
      1 svartaktig
      5 svartbrun
      2 svartbrunt
      1 svartfärgad
      1 svartglansigt
      1 svartgrön
      1 svårtillgänglig
      1 svartkroppsstrålning
      1 svartlut
      1 svartmagi
      1 svartmarkerade
      1 svartnade
      1 svärtning
      1 svårtolkad
      2 svartpest
      1 svartpolerat
      2 svartråttan
      5 svartsjuka
      2 svartsjukan
      1 svartsjuke
      1 svartsoppa
      1 svartvattenfeber
      2 svartvioletta
      1 svartvit
      1 svartvita
      1 svartvitt
      1 svårundersökt
      1 svårutredd
      1 svårutrotad
      1 svåruttalade
      1 svarvad
      1 svarvning
      1 svävande
      3 svävar
      7 svavel
      1 svavelatomen
      1 svavelatomer
      1 svavelbindningar
     13 svaveldioxid
      1 svaveldioxidens
      1 svaveldioxidmolekylen
      1 svaveldioxidutsläppen
      1 svavelfattig
      1 svavelföreningar
      1 svavelgul
      4 svavelhaltiga
     19 svavelsyra
      1 svavelsyran
      1 svavelsyrebindningen
      1 svavelsyrlighet
      1 svaveltillsatsen
      2 svaveltrioxid
      4 svavelväte
      1 svbk
      1 svd
      1 sve
      1 svealands
      1 sveavägen
     10 sveda
      1 sveen
      2 sven
      1 sveninge
      1 svenner
      1 svenolov
      1 svenshögens
     83 svensk
    265 svenska
      9 svenskan
      3 svenskans
     17 svenskar
      3 svenskarna
      1 svenskbrittisk
      1 svenskdanske
     11 svenske
      4 svensken
      1 svenskneurootologiskförening
      2 svenskspråkiga
      9 svenskt
      1 svep
      1 svepavstämda
      1 svepe
      1 svepeblad
      1 svepen
      1 sveper
      1 svepet
      1 svepets
      1 svepgenerator
      1 svephastigheten
      1 sveps
      3 svepte
      1 sverak
    984 sverige
      1 sverigeref
     65 sveriges
      3 sves
      1 svetsade
      1 svetsas
      2 svetsning
     29 svett
      1 svettämnen
     10 svettas
      1 svettdrivande
      1 svetteduk
      4 svetten
      1 svettens
      1 svettig
      1 svettkanalerna
      1 svettkörtelns
     10 svettkörtlar
      2 svettkörtlarna
      1 svettlukten
      2 svettmängd
      2 svettmängden
      1 svettmängder
     21 svettning
     19 svettningar
      2 svettningen
      1 svettutsöndring
      1 svettvätskan
      1 svida
      2 svider
      2 svikit
      1 svikt
      1 svikta
      3 sviktande
      2 sviktar
      1 svimfärdig
      4 svimma
      1 svimmade
      1 svimmande
      5 svimmar
     11 svimning
      3 svimningar
      1 svimningarna
      6 svin
      1 svinbandmask
      2 svindel
      1 svindla
      1 svindlande
      1 svinga
      2 svinhår
      5 svininfluensa
      1 svininfluensaepidemin
      2 svininfluensan
      4 svinkoppor
      1 svinmålla
      1 sviter
      2 sviterna
      1 svkomododrake
      1 svordomar
      2 svt
      5 svullen
      1 svullet
     25 svullna
     53 svullnad
      2 svullnade
     18 svullnaden
      4 svullnader
      1 svullnaderna
     12 svullnar
      1 svullnartäpps
      6 svulst
      1 svulstartade
      1 svulstcellerna
      2 svulsten
      2 svulsterna
      1 svulstfall
      1 swäfande
      2 swahili
      1 swahiliska
      6 swami
      1 swåra
      1 swarfarin
      1 swaziland
      1 sweden
      1 swedenborg
      1 swedish
      1 swedo
      1 sweep
      2 swift
      1 swisnfkomplexet
      1 swiss
      3 sy
      6 sycosis
      7 syd
      9 sydafrika
      1 sydafrikanågra
      2 sydafrikanska
     23 sydamerika
      2 sydasien
      1 sydcentrala
      1 sydda
      1 syddansk
      2 sydde
      5 sydenham
      2 sydenhams
      1 sydeuropa
      1 sydeuropéerna
      1 sydeuropeiska
      2 sydgullregn
      1 sydgullregnets
      5 sydkorea
      1 sydkoreanska
      1 sydlig
      2 sydliga
      3 sydligaste
      1 sydney
      1 sydöst
      1 sydostasiater
      9 sydostasien
      1 sydostasiens
     11 sydöstra
      1 sydpolen
      1 sydsec
      1 sydspets
      1 sydssverige
      1 sydsvenska
      1 sydsverige
      2 sydtyrolens
      7 sydvästra
     97 syfilis
      2 syfilisbakterier
      1 syfilisbehandling
      3 syfilisen
      1 syfilisepidemi
      1 syfilisexperiment
      1 syfilisgener
      1 syfilisinfektion
      1 syfilisproteiner
      1 syfilissåret
      1 syfilissmitta
      2 syfilissmittade
      1 syfilistester
      3 syfilitisk
      1 syfilitiska
     17 syfta
      6 syftade
      3 syftande
    108 syftar
     91 syfte
     10 syften
      1 syftena
     41 syftet
      2 syftning
      1 sykehus
      1 sykepleie
      1 sylar
      2 sylt
      1 sylvain
      1 sylvania
      1 sylvaticum
      1 sylvestris
      1 sylvia
      1 symaskinen
      2 symbionter
      2 symbios
      1 symbiotiska
      1 symbiotiskt
     16 symbol
      6 symbolen
     11 symboler
      6 symbolerna
      1 symbolik
      1 symboliken
      2 symboliserade
      1 symboliserar
      1 symboliseras
      1 symboliserats
      2 symbolisk
      4 symboliska
      2 symbolspråk
      1 symbolspråken
      1 symfonier
      1 symfoniorkester
      1 symfoniorkesters
      1 symfysen
      1 symfyseolys
      1 symfyseolyslesioner
      2 symfyseotomi
      1 symfyseotomin
      1 symfysis
      3 symmetrisk
      1 symmetriska
      1 symmetriskt
      2 sympati
      1 sympaticuspåslag
      1 sympatikuspåslag
     14 sympatiska
      1 symphysis
      1 symposier
      1 symposion
    447 symptom
      1 symptomatisk
      3 symptomatiska
      1 symptombeskrivningen
      2 symptombild
      5 symptombilden
      1 symptombilder
      2 symptomdebut
    169 symptomen
      3 symptomens
     24 symptomet
      5 symptomfri
      5 symptomfria
      1 symptomfrihet
      3 symptomfritt
      1 symptominriktad
      2 symptomlindrande
      1 symptomlindring
      1 symptomlös
      1 symptomreduktion
      1 symptomtetraden
      1 symptomutslaget
      1 sympton
    421 symtom
      8 symtomatisk
     10 symtomatiska
      3 symtomatiskt
      1 symtomatologin
      7 symtombild
      2 symtombilden
      1 symtombilder
      4 symtomdebut
      1 symtomdefinitioner
    154 symtomen
      4 symtomens
      1 symtomer
     12 symtomet
      5 symtomfri
      7 symtomfria
      1 symtomfrihet
      4 symtomgivande
      1 symtomlindrande
      1 symtomlindrare
      2 symtomlindring
      1 symtomlös
      1 symtomreducering
      1 symtomreduktion
     63 syn
      7 synanon
      1 synanonmedlemmar
      1 synapomorfi
      8 synaps
      3 synapsen
     14 synapser
      1 synapserna
      1 synapsgapet
      1 synapsklyfta
      4 synapsklyftan
      1 synapskopplingar
      1 synapsplasticiteten
      1 synapsspalten
      1 synapsspatiet
      1 synapsspringan
      1 synaptisk
      5 synaptiska
      4 synas
      2 synbar
      3 synbara
      1 synbarligen
      1 synbart
      1 synbesvär
      1 synbeteende
      3 synbortfall
      1 syncellerna
      1 syncentralerna
      1 syncope
      3 syncytialvirus
      1 syncytialviruset
      1 synd
      1 syndactyli
      3 syndaktyli
      1 syndat
      2 synder
      2 synderna
      1 syndig
      1 syndigt
    199 syndrom
     18 syndrome
      1 syndromen
      4 syndromes
     29 syndromet
      2 syndromets
      1 syndromklassificering
     30 synen
      1 synergieffekt
      1 synergieffekter
      1 synergonomiska
      5 synes
      2 synestesi
     11 synfält
      1 synfälten
     13 synfältet
      2 synfältsbortfall
     12 synfel
      1 synfelet
      1 synförändringar
      1 synförlust
      2 synförmåga
      1 synförsämring
      1 synfunktion
      1 syngami
      1 synhallucination
      7 synhallucinationer
      1 synhallucinationerna
      4 synhjälpmedel
      6 synintryck
      1 synintrycken
      1 synkomfort
      3 synkope
      1 synkopering
      1 synkron
      1 synkronisera
      1 synkroniserade
      1 synkroniserar
      1 synkronisering
      2 synkrotron
      8 synlig
     20 synliga
      1 synliggör
      1 synliggöra
      1 synliggöras
      1 synliggörs
      4 synligt
      7 synnedsättning
     98 synnerhet
      1 synnerlig
      7 synnerligen
      1 synnerv
      3 synnerven
      1 synnervens
      1 synnervsinflammation
      1 synnervskorset
      1 synomfånget
     17 synonym
      1 synonyma
     22 synonymer
      1 synonymis
     27 synonymt
      1 synoskärpa
      1 synpåverkan
      3 synproblem
      6 synpunkt
      1 synrester
      3 synrubbningar
     47 syns
     22 synsätt
      1 synsätten
      9 synsättet
      1 synsinnet
      5 synskada
      1 synskadad
      1 synskadadade
      5 synskadade
      4 synskadades
      8 synskärpa
      6 synskärpan
      1 synskärpeavståndet
      2 synstörningar
      1 synsymptom
      1 syntaxordföljd
     16 syntes
     20 syntesen
      1 syntesgas
      1 synteshastigheten
      1 syntesråvara
      1 syntester
      2 syntesväg
      1 syntet
      1 syntetborste
      1 syntetfiber
      3 syntetisera
      1 syntetiserade
      3 syntetiserades
      3 syntetiserar
     10 syntetiseras
      1 syntetiserats
      1 syntetisering
      1 syntetiseringen
      1 syntetisk
     18 syntetiska
     16 syntetiskt
      1 syntetmaterial
      1 syntton
      6 synvinkel
      1 synvinkeln
      1 syphilis
      1 syphilus
      9 syra
      1 syraangrepp
      1 syraattacker
      1 syrabasbalans
      1 syrabasbalansen
      1 syrabasbalasen
      1 syrabasrelationen
      1 syrabehandling
      1 syrade
      2 syrafast
      3 syrafasta
      1 syraförgiftning
      1 syraform
      1 syrahämmande
      1 syrakänsliga
      1 syrakatalyserad
      1 syraklorider
      1 syrakoncentrationen
      2 syrakonstant
      1 syrakonstanten
      1 syramantel
      9 syran
      1 syrans
      1 syras
      1 syrasekretionshämmarna
     87 syre
      2 syreatom
      2 syreatomer
      1 syrebärare
      1 syrebaserade
      2 syrebehov
      1 syreberikad
     28 syrebrist
      1 syrebristen
      5 syrefattig
      5 syrefattiga
      6 syrefattigt
      1 syreförbrukning
      1 syrefri
      1 syrefrisättning
      1 syrehalt
      3 syrehalten
      2 syrehemoglobindissociationskurvan
      3 syrekoncentrationen
      1 syreluft
      1 syremättnad
      2 syremättnaden
      1 syremättnadsgrad
      1 syremolekyl
      1 syrenivå
      2 syrenivån
      1 syreomsättningen
      2 syreradikalerna
      1 syrerik
      3 syrerika
      4 syrerikt
      2 syresatt
      2 syresatta
      8 syresätta
      2 syresätter
      7 syresättning
      3 syresättningen
      1 syresatts
      3 syresätts
     11 syret
      3 syretillförsel
      1 syretransport
      1 syretransporten
      1 syretransporterande
      1 syretryck
      2 syretrycket
      4 syrets
      1 syreupptag
      1 syreupptaget
      3 syreupptagningsförmåga
      2 syreupptagningsförmågan
      1 syreutvinning
     55 syrgas
      1 syrgasbehandling
      2 syrgasbrist
      1 syrgasens
      3 syrgasförgiftning
      1 syrgasgrimma
      2 syrgashalt
      1 syrgashalten
      1 syrgaskoncentration
      1 syrgaskoncentrationen
      5 syrgasmättnad
      1 syrgasmättnaden
      2 syrgasmolekyl
      2 syrgasmolekylen
      3 syrgasmolekyler
      1 syrgasnivåer
      1 syrgaspartialtrycket
      1 syrgassensor
      2 syrgastransport
      1 syrgastransporten
      2 syrgasupptag
      4 syrien
      2 syringomyeli
      1 syringomyelia
      1 syriska
      1 syrlig
     14 syror
      7 sys
     11 syskon
      1 syskonspråkens
      1 sysselsätta
      1 sysselsatte
      7 sysselsättning
      1 sysselsättningar
      1 sysselsättningsterapi
      1 sysselsätts
      1 syssla
      2 sysslade
      8 sysslar
      1 sysslolös
      4 sysslor
     90 system
      2 systema
      1 systematic
      6 systematik
      1 systematisera
      1 systematiserade
     16 systematisk
     13 systematiska
     24 systematiskt
      1 systembolaget
      1 systemcirkulationen
      5 systemen
     65 systemet
      1 systemets
      1 systemfelen
      9 systemisk
      9 systemiska
      2 systemiskt
      6 systemkretsloppet
      1 systemkretsloppetvar
      2 systems
      3 syster
      1 systerklass
      1 systertaxon
      1 systole
      1 systolefasen
      1 systoliska
      1 sytomerna
      4 szasz
    145 t
      1 [t]
    338 ta
      1 tá
     13 tå
      1 tabacum
      1 tabakobon
      3 tabell
      3 tabellen
      1 tabernanthe
      2 tabes
     13 tablett
      5 tabletten
     26 tabletter
      6 tabletterna
      6 tablettform
      2 tablettintag
      1 tablettintaget
      1 tablettmaskin
      1 tablettöverdos
      1 tabloiden
      5 tabu
      2 tabubelagd
      2 tabubelagt
      4 tabun
      1 tabut
      1 tac
     35 tack
     10 täcka
      1 tackan
      2 täckande
      1 täckas
      1 tacke
      1 täcken
     26 täcker
      1 täckmantel
      1 täckning
      3 tackor
     11 täcks
      1 tacksamma
     12 täckt
      8 täckta
      3 täckte
      1 tacos
      1 tadeusz
      1 tado
      1 taekwondo
      2 taenia
      1 taföreningen
      1 taft
     29 tag
     10 tåg
      1 tagande
      3 tagen
      1 tages
     33 taget
      7 tåget
      1 tagetes
      3 tågets
      5 taggar
      1 taggig
      1 taggiga
     47 tagit
     20 tagits
      1 tagliacozzi
      2 tagna
      1 tagning
      2 tågolyckor
      1 tågresor
      1 tågtrafik
      2 tai
      1 taigafästing
      1 taipan
      4 taipanen
      2 taipaner
      3 taiwan
      8 tak
      1 taken
      5 taket
      2 takfallet
      1 takk
      1 takläggare
      1 taklyftar
      1 takman
     35 takt
      1 taktäckning
      1 taktäckningsändamål
      1 taktegellika
      2 taktik
      1 taktiken
      1 taktiker
      4 taktil
      4 taktila
      1 taktilt
      1 taktisk
      3 taktiska
      1 taktslag
      7 takykardi
      4 takypné
    116 tal
     20 tål
     22 tala
      7 tåla
      1 talad
     10 talade
      1 talamisk
      2 tålamod
     33 talamus
      4 talande
      1 talapparat
      4 talapparaten
      1 talapparatens
      3 talapraxi
     71 talar
      3 talare
      1 talaren
      1 talarens
      1 talares
      7 talas
      1 tålas
      6 talassemi
      1 �talassemi
      2 talassemier
      6 talat
      3 talböcker
      1 talbok
      1 talboken
      3 talboks
      1 talcum
      1 tåleder
     17 talen
      1 �talen
      1 talesättet
      1 talessätt
      1 talessemi
    750 talet
      1 talét
     33 talets
      1 talflöde
      1 talflödet
      1 talförbättrande
      1 talförmåga
      1 talförståelse
      4 talg
      1 talgestaltare
      7 talgkörtlar
      2 talgkörtlarna
      2 talhandling
      1 taliaferro
     24 talidomid
      3 tålig
      1 tålighet
      3 tåligt
      1 talionprincipen
      1 talisterna
      4 täljsten
     12 talk
      1 talkaraktär
      1 talkbox
      2 talkpuder
      3 tall
      1 talläten
      1 tallbarr
      2 talljud
      1 talljudet
      1 tallkärneolja
      5 tallkottkörteln
      1 tallkottskörtel
      2 tallrikar
      1 tallriken
      1 tålmodiga
      1 talmotoriken
      1 talmuskler
      2 talorgan
      2 talorganen
      1 talorganens
      1 talpedagog
      2 talproduktion
      1 talproduktionen
      4 talrädsla
      1 talrik
      3 talrika
      3 talröret
      1 talrörsestimering
      2 talröst
      1 talrytm
      1 talrytmstörningar
      2 tals
      1 talserien
      1 talsfilmer
      1 talsfilosofen
      1 talsforskare
      2 talsfysiologen
      2 talshus
      1 talsituationen
      5 talspråk
      2 talspråket
      1 talspråkliga
      3 talstörning
      2 talstörningar
      1 talsutgåvans
      6 talsvårigheter
      1 talsvårigheterna
      1 talsyntes
      1 talsyntesprogram
      1 tält
      2 talteknologi
      1 talterapeut
      1 talträningsändamål
      1 talutveckling
      1 tama
      1 tamar
      1 tamaulipa
      1 tambin
      4 tamboskap
      3 tamdjur
      1 tåmellanrum
      2 tamfår
      1 tamgris
      1 tamgrisen
      1 tamhundar
      2 tamiflu
     34 tämligen
      1 tammi
      2 tamoxifen
      1 tamponad
      8 tampong
      2 tamponganvändning
      6 tampongen
     15 tamponger
      1 tampongludd
      1 tampongsjukan
      1 tamsvin
      1 tamt
      5 tån
      1 tanach
      1 tånaglar
      1 tånaglarna
      3 tand
      8 tända
      3 tandade
      1 tändande
      1 tandanlag
      1 tandarbete
      1 tändare
      1 tandbehandlingar
      1 tandbehandlingsmaterial
      1 tandbenet
      1 tandbettet
      8 tandblekning
      1 tandblekningsmedel
      1 tandblekningsmetoder
      1 tandblekningspenna
      1 tandblekningsprodukter
      1 tandborr
      4 tandborstar
     12 tandborste
      9 tandborsten
      1 tandborstens
      1 tandborsthuvudet
     12 tandborstning
      2 tandborstningen
      1 tandbryggor
      1 tandemaljen
      1 tandemaljprover
      6 tanden
      1 tandens
     60 tänder
      1 tänderkäkar
     83 tänderna
      6 tändernas
      1 tandersättningar
      1 tandfästet
      1 tandfickorna
      1 tandförlust
      2 tandfyllningar
      3 tandgnissling
      1 tandhälsan
      2 tandhalsar
      1 tandhälsoinformation
      1 tandhalsytan
      1 tändhatt
      2 tandhygien
      9 tandhygienist
      1 tandhygienisten
      1 tandhygienister
      1 tandhygienistyrket
      1 tandimplantat
      1 tandinfektioner
      1 tandkaries
      1 tandkarpar
      1 tandkitt
      8 tandkött
     13 tandköttet
      1 tandköttets
      1 tandkötts
      1 tandköttsfickor
      4 tandköttsinflammation
      1 tandköttsinflammationer
      1 tandköttsirritation
      2 tandköttskanten
      1 tandköttsproblem
     32 tandkräm
      6 tandkrämen
      6 tandkrämer
      1 tandkronor
      2 tandlagningar
      1 tandlagningsamalgam
      4 tandläkarbesök
      2 tandläkarborren
      1 tandläkarbrist
     49 tandläkare
      9 tandläkaren
      2 tandläkarens
      3 tandläkarexamen
      3 tandläkarförbund
      1 tandläkarförbunds
      1 tandläkarinstrument
      1 tandläkarkåren
      1 tandläkarkunskap
      2 tandläkarlegitimation
      2 tandläkarna
      1 tandläkarnas
      4 tandläkarskräck
      1 tandläkarstudenter
      2 tandläkarutbildning
      3 tandläkarutbildningen
      1 tandläkarvetenskap
      4 tandläkaryrket
     12 tandlossning
      1 tandlossningssjukdom
      1 tandlossningssjukdomarna
      1 tandmasken
      1 tandmellanrum
      1 tändningsläget
      1 tandnyckel
      1 tandömsning
      1 tandpasta
      2 tandpetare
      1 tandplack
      1 tandpressning
      1 tandprotes
      1 tandproteser
      1 tandpulver
      1 tandrad
      1 tandraden
      1 tandreglerande
      2 tandreglerare
      3 tandreglering
      3 tandregleringen
      1 tandröntgenundersökning
      2 tandröta
      1 tandsällning
      1 tandsjukdomar
      2 tandskena
      3 tandsköterska
      3 tandsköterskan
      1 tandsköterskeutbildningar
      1 tandsköterskor
      1 tandskydd
      1 tandskyddet
      1 tandsmärtorskador
      7 tandställning
      5 tandställningar
      9 tandställningen
      1 tandstatus
     12 tandsten
      2 tandstenen
      4 tandsticka
      3 tändsticka
      1 tandstickan
      1 tandstickor
      1 tändstickorna
      2 tändsticksaskar
      1 tändsticksaskarna
      1 tandsubstans
      1 tandsubstansen
      2 tandtekniker
      1 tandteknisk
     17 tandtråd
      4 tandtråden
      1 tandtrådshållare
      1 tandupplysningen
     17 tandvård
      7 tandvården
      3 tandvårdens
      1 tandvårds
      1 tandvårdsfobi
      1 tandvårdsinstitutet
      1 tandvårdskostnader
      2 tandvårdsrädsla
      4 tandvärk
      1 tandvärkstallar
      1 tandytan
      1 tandytorna
      3 tång
      4 tångamperemeter
      3 tångamperemetern
      2 tångamperemetrar
      1 tångaska
      2 tången
      1 tångens
      1 tangerade
      1 tangerar
      1 tånghalvor
      1 tångliknande
      1 tångskaften
      1 tänja
      2 tänjer
      1 tänjning
      6 tänjs
      1 tänjt
      2 tank
      3 tänk
     35 tänka
     25 tänkande
      1 tänkanden
      5 tänkandet
     85 tankar
      3 tänkare
     18 tankarna
      4 tänkas
      2 tänkbar
      6 tänkbara
      1 tänkbart
     20 tanke
      1 tankebanorna
      1 tankeblockering
      3 tankedetraktion
      1 tankeeko
      1 tankefältterapi
      6 tankeflykt
      1 tankeförloppsstörning
      2 tankeförmåga
      3 tankeförmågan
      1 tankefunktion
      1 tankegångar
      1 tankegångarna
      1 tankegången
      2 tankeinnehåll
      2 tankeliv
      6 tankelivet
      1 tankemönstren
     25 tanken
      3 tankepåsättning
      1 tankeprocesser
      1 tankeprocesstörning
     14 tänker
      1 tänkes
      3 tankesätt
      1 tankesättet
      2 tankestopp
      7 tankestörning
     21 tankestörningar
      1 tankestörningarna
      1 tanketråden
      1 tanketröghet
      1 tankeutbredning
      1 tankevärld
      2 tankeverksamhet
      1 tankeverksamheten
      1 tanklig
      1 tanklöshet
      1 tankmetoden
      2 tänks
     13 tänkt
      3 tänkta
      2 tänkte
      1 tanlines
      2 tanner
      4 tannerskalan
      1 tänt
      1 tantrisk
      1 tantriska
      1 tantriskt
      7 tanzania
      1 tao
      1 taorganisation
      1 tapas
      1 tapet
      1 taphrina
      1 tapp
     11 tappa
      6 täppa
      2 tappade
      2 tappades
     16 tappar
      3 tappas
      3 täppas
      6 tappat
      2 tappats
      3 tappen
      4 täpper
      2 tappning
      1 tappningar
      3 tappningen
      1 tappningkatetrarna
      1 tappningsaggregatet
      1 tappningskateter
      3 tappningskatetrar
      1 tappningspåsen
      5 täpps
      1 tappstället
      2 täppt
      1 täppts
    303 tar
     18 tår
      1 tära
      2 tarandi
      1 tarantel
      2 tarantella
      1 tarantism
      1 tarantismen
      1 taranto
      1 tarantula
      1 tårar
      1 tardigrader
      3 tardiv
      1 tardiva
      1 tårflöde
      1 tårgas
      1 targeted
      2 targets
      1 tarjei
     19 tarm
     10 tarmar
     22 tarmarna
      1 tarmarnas
      2 tarmavsnitt
      6 tarmbakterier
      4 tarmcancer
      1 tarmceller
      2 tarmdel
      1 tarmdelen
     90 tarmen
     17 tarmens
      1 tarmfickor
      7 tarmflora
     14 tarmfloran
      9 tarmflorans
      1 tarmförträngningar
      1 tarmfunktion
      1 tarmfunktionen
      1 tarmfunktioner
      1 tarmhåligheten
      2 tarminfektion
      1 tarminfektioner
      4 tarminflammation
      3 tarminnehåll
      9 tarminnehållet
      2 tarminnehållets
      3 tarmkanal
     28 tarmkanalen
      3 tarmkanalens
      1 tarmkäx
      4 tarmkäxet
      1 tarmkirurgi
      1 tarmkrökarna
      1 tarmloppet
      2 tarmludd
      2 tarmlumen
      1 tarmlymfa
      1 tarmmotorik
      1 tarmopererade
      1 tarmöppningen
      1 tarmparasit
      1 tarmplack
      3 tarmproblem
      6 tarmrening
      1 tarmresektioner
      1 tarmretande
      1 tarmrörelser
      5 tarmrörelserna
      9 tarmsjukdom
      7 tarmsjukdomar
      1 tarmsköljningar
      1 tarmsköljningsmedel
      2 tarmslemhinna
      2 tarmslemhinnan
      3 tarmslemhinnans
      1 tarmslemmhinor
      1 tarmslingan
      2 tarmstopp
      2 tarmsuturer
      1 tarmsuturerna
      3 tarmsvikt
      1 tarmsymtom
     14 tarmsystemet
      7 tarmtömning
      1 tarmtrådars
      1 tarmtuberkulos
      1 tarmvägg
      2 tarmväggarna
      9 tarmväggen
      1 tarmväggens
      1 tarmvätskan
      1 tarmvilli
      6 tarmvred
     13 tårna
      1 tarnier
      1 tarniers
      1 tärningar
      1 tärnsjö
      1 tårs
      1 tårsubstitut
      1 tärt
      1 tårvätskan
    169 tas
      1 task
      1 tåskador
      1 tasmanske
      1 tassen
      1 tassinlademilune
      6 tät
     14 täta
      1 tätar
      5 tätare
      1 tätbefolkat
      4 täthet
      1 täthetskillnaderna
      1 tåtila
      1 tätnar
      1 tätning
      1 tätort
      1 tätorter
      1 tätslutande
      1 tatsurou
     36 tätt
      1 tattare
      1 tattoe
      1 tattoo
      1 tättslutande
      3 tatuera
      4 tatuerare
      1 tatuerares
      9 tatuering
      5 tatueringar
      2 tatueringen
      1 tatueringsfärg
      1 tatueringsfärgeninket
      1 tatueringsfärger
      1 tatueringsstudior
      2 tatueringstillfället
      2 tatula
      1 tätvuxna
      1 taupin
      1 tauricola
      1 taurin
      1 tautomeriska
      1 tavelformade
      2 tavistockkliniken
      1 tävla
      1 tävlar
      1 tävlare
      1 tävlas
      1 tävlat
      5 tävling
      3 tävlingar
      1 tävlingsgrenar
      1 tävlingsinriktade
      1 tävlingsinstinkt
      1 tävlingsperiod
      2 tavlor
      1 taxaner
      1 taxering
      1 taxichaufförers
      1 taxin
      2 taxol
      1 taxonomi
      1 taxonomiskt
      1 taxonomy
      4 taxus
      2 tb
      4 tbc
      8 tbe
      1 tbefall
      1 tbeföreningen
      1 tbeinfektion
      2 tbesmitta
      1 tbesmittade
      3 tbg
     11 tbt
      1 tbtbemålat
      1 tbtrelaterade
      1 tc
      4 tca
      1 tcaantidepressiva
     11 tceller
      1 tcellerml
      3 tcellerna
      1 tcells
      1 tcellslymfom
      1 tcfl
      1 tchadsjön
      1 tcm
      1 tco
      1 tcomärkning
      1 tcos
      1 tcotidningen
      2 tdd
      1 tddelektroder
     11 te
      3 teaching
     14 team
      1 teamen
      1 teamens
      4 teamet
      1 teammodell
      2 teater
      1 teatern
      1 teaterpjäs
      1 teaterroller
      1 teatersmink
      1 teatraliskt
      1 teatrar
      1 tebain
      1 tebuskens
      1 teceremonin
      1 tech
      1 technegas
      1 technical
      1 technologies
      1 technos
    175 tecken
      1 teckenet
      8 teckenspråk
      1 teckenspråket
      2 teckenspråkiga
      3 tecknad
      1 tecknade
      1 tecknande
      1 tecknar
      2 tecknas
      2 tecknat
     12 tecknen
     11 tecknet
      1 teckning
      5 teckningar
      1 teckningen
      1 ted
      3 tee
      1 teflon
      2 teg
      2 tegel
      1 tegelsten
      2 tegenero
      1 tegmentområdet
      1 teichoic
      1 teicoplanin
      2 tein
      1 tej
      2 tejp
      1 tejpa
      1 tejpar
      1 tejpas
      1 tejpbit
      1 tejpen
      1 tejpprov
      1 tekken
      7 teknetium
      2 teknetiumm
      1 teknetiummgeneratorer
      1 teknetiumviisukfid
     65 teknik
     28 tekniken
      2 teknikens
     28 tekniker
      1 teknikern
      2 teknikerna
      1 tekniknivå
      1 teknikorienterade
      1 teknikstress
     18 teknisk
     19 tekniska
      1 tekniskaarbetshygieniska
     11 tekniskt
      3 teknologi
      2 teknologin
      1 tekom
      1 tekopp
      1 tekoppar
      1 tektonisk
      3 tektronix
      1 tele
      7 telefon
      1 telefonanalysprogram
      2 telefoner
      1 telefonjourer
      1 telefonkommunikation
      1 telefonkontakt
      1 telefonkvalitet
      1 telefonlinjer
      1 telefonlur
      1 telefonlurar
      1 telefonnummer
      1 telefonrådgivande
      1 telefonrådgivning
      1 telefonsamtal
      1 telefonsamtalsregister
      2 telefonstöd
      1 telefonstödet
      1 telegrafister
      3 telehälsa
      1 teleknetiska
      1 telekomindustrin
      1 telekommunikationsföretag
      1 telekommunikationsutrustning
      1 telemark
      6 telemedicin
      1 telepatisk
      1 telepatiska
      1 telepatiskt
      1 teleskopord
      1 teleslingor
      1 telespole
      1 televerket
      4 tema
      9 teman
      1 temat
      1 tematiskt
      1 temgesic
      1 temomätning
      1 tempeh
      7 tempel
      1 tempelbyggnader
      1 tempeldanser
      1 tempellivet
      3 temperament
      1 temperamentet
     49 temperatur
      2 temperaturbaserade
      1 temperaturberoende
      1 temperaturcentrum
      1 temperaturchocker
     16 temperaturen
     24 temperaturer
      1 temperaturerna
      1 temperaturförändringar
      1 temperaturinställningar
      1 temperaturisolerande
      1 temperaturkänsligheten
      1 temperaturökningen
      1 temperaturreglering
      1 temperaturregleringen
      1 temperatursänkning
      1 temperaturstegring
      1 temperaturvariationer
      1 temperaturväxlingar
      5 tempererade
      3 tempererat
      3 templat
      1 templatet
      2 templet
      9 tempo
      2 temporal
      1 temporalis
      2 temporalloben
      1 temporallobennedre
      3 temporalloberna
      2 temporallobsepilepsi
      1 temporallobsresektion
      6 temporär
      1 temporära
      6 temporärt
      2 tempot
     20 tendens
      2 tendensen
      1 tendenser
      1 tendenserna
      2 tenderade
     40 tenderar
      1 tenderat
      2 tenn
      1 tennatom
      2 tennessee
      1 tennfluorid
      1 tennföreningar
      1 tennis
      1 tennisarm
     14 tennisarmbåge
      1 tennisplan
      1 tennisracket
      1 tennisracketar
      1 tennisracketen
      2 tennisspel
      1 tennisspelares
      1 tennjon
      9 tens
      1 tensapparat
      2 tensider
      1 tension
      1 tenssmärtlindring
      1 tentakel
      1 tentakellängden
      5 tentakler
      4 tentaklerna
      2 tentamen
      1 tentativt
      1 tenue
     13 teobromin
      1 teobrominet
      3 teobrominförgiftning
      1 teodicé
      1 teodolitgoniometrar
      1 teofyllaminpreparat
      1 teofyllin
      3 teologer
      3 teologi
      2 teologin
      2 teologisk
      1 teologiska
      1 teologiskt
      2 teoretiserande
      1 teoretiserat
      1 teoretiserats
      6 teoretisk
      9 teoretiska
     10 teoretiskt
     62 teori
      2 teoribildning
      1 teoribildningen
     42 teorier
      8 teorierna
     46 teorin
      1 teorins
      1 teos
      1 teosofin
      1 teosofins
      1 tephrosia
      2 tequila
      1 tequilaagave
      1 tequilana
      4 ter
      1 tera
      1 terapand
      3 terapeut
     11 terapeuten
      4 terapeutens
      3 terapeuter
      1 terapeuterna
      8 terapeutisk
     11 terapeutiska
      3 terapeutiskt
     49 terapi
      7 terapier
      8 terapiform
      3 terapiformen
      6 terapiformer
      1 terapiformerna
      1 terapiforskning
      6 terapihund
      1 terapihundar
      3 terapihunden
      2 terapimetod
     17 terapin
      1 terapiresistenta
      1 terapisessioner
      1 terapiverksamhet
      2 teras
      1 teratogena
      2 teratogener
      1 teratogenicitet
      2 teratologi
      7 teratom
      1 terence
      1 teresa
      4 teriak
     57 term
    108 termen
      1 termens
     26 termer
     10 termerna
      1 termin
      3 terminal
      3 terminala
      1 terminalen
      2 terminalt
      5 terminer
     14 terminologi
      1 terminologimässigt
      5 terminologin
      1 terminologiråd
      3 termisk
      3 termiska
      1 termiskt
      1 termodynamikens
      1 termodynamiska
      1 termogenin
      1 termohypestesi
      1 termokauterisering
      1 termokoagulation
      1 termoplast
      1 termoplegi
      1 termoreceptorer
      1 termoreceptorerna
      3 termoreglering
      5 termoregleringen
      2 termostat
      1 termostatreglerade
      1 termostatstrykjärnet
      1 terpen
      1 terpentin
      1 terrakotta
      1 terramycin
      1 terrängen
      1 terrarium
      1 terre
      2 territorier
      3 territorium
      1 territory
      1 terror
      1 terrorattacker
      1 terroriserade
      1 terrorism
      1 terroristbekämpningen
      1 terrorister
      1 terrorn
      2 ters
      1 tertbutanol
      5 tertiär
      6 tertiära
      1 tertiärförebyggande
      2 tertiärt
      1 terveyskeskus
      2 tes
      3 tesen
      1 teser
      1 tesked
      1 tesorten
     83 test
     11 testa
      5 testade
      6 testades
      1 testamente
     10 testamentet
      1 testamentets
      4 testar
     22 testas
      2 testat
     13 testats
      1 testbildsgeneratorn
      1 testdata
      8 testen
     48 tester
      7 testerna
      1 testernas
     27 testet
      4 testikel
      1 testikelcancer
      4 testikelinflammation
     19 testikeln
      2 testikelns
      1 testikeltorsion
      1 testikeltumör
      1 testikelvävnaden
     16 testiklar
     46 testiklarna
      4 testiklarnas
      1 testis
      1 testisretention
      4 testistorsion
      1 testmedicinen
      2 testmetod
      1 testmetoden
      3 testmetoder
      1 testmetods
      4 testning
      1 testningen
     88 testosteron
      1 testosteronaktiviteten
      1 testosteronbaserade
     12 testosteronbrist
      1 testosteronbristen
     14 testosteronet
      7 testosteronets
      1 testosteronhalt
      1 testosteronindex
     12 testosteronnivåer
      5 testosteronnivåerna
      1 testosteronnviåer
      1 testosteronpreparat
      1 testosteronproduktionen
      1 testosteronreceptorn
      1 testosteronreglering
      1 testosteronresistens
      1 testosterontillförsel
      3 testosteronvärden
      1 testpanel
      4 testpersonen
      1 testpersoner
      1 testpersons
      7 testresultat
      1 testresultaten
      1 teststickor
      1 teststickorself
      1 testterminologin
      1 testurval
      1 tesvamp
      1 tet
      4 tetani
      2 tetanus
      2 tetanustoxin
      2 tetanustoxinet
      1 tetra
     10 tetracyklin
     12 tetracykliner
      1 tetracyklinerev
      1 tetracyklinerna
      1 tetracyklinresistens
      1 tetradehydro�epoximetoximetylmorfinanol
      1 tetraetylbly
      1 tetrafluoretan
      2 tetrafluoreten
      1 tetragonalt
      1 tetrahydrobiopterin
      1 tetrahydrofolat
      1 tetrakloretan
      1 tetraklormetan
      1 tetralin
      1 tetramer
      1 tetraoxidifenylmetankarboxylsyra
      1 tetraplegi
      1 tetraplegiker
      1 tetrapyrrol
      2 tetrapyrroler
      1 tetrapyrrolsyntesen
      1 tetrasomi
      2 tetrasomier
      1 tewtraining
    120 tex
      5 texas
     10 text
      1 textböcker
     13 texten
      9 texter
      3 texterna
      1 textfunktionsmjukvara
      2 textil
      1 textilfärgning
      1 textilhanddukar
     22 textilier
      2 textilierna
      1 textilindustrin
      1 textilis
      1 textilt
      1 textiltvätt
      1 textiltypen
      1 textilvara
      1 textkanon
      1 textpartier
      1 texttelefon
      1 texttelefoner
      1 texttelefoni
      1 texttelefonsamtal
      1 texturer
      1 tfpi
      1 tft
      2 tg
      1 tgak
      1 tgf
      1 tgn
      1 thai
      8 thailand
      1 thailändska
      4 thalamus
      1 thalamusfunktion
      1 thalamuskärnor
      1 thalassa
      2 thalassemi
      2 thalidomid
      1 than
      7 that
      1 thc
      1 thdominerad
    126 the
      2 theca
      1 thecacellerna
      1 their
      1 thell
      1 thelpercells
      1 them
      1 themsen
      2 theodor
      1 théophile
      1 theophrastus
      1 theorein
      2 theory
      1 theralen
      2 therapeia
      1 theraphy
      1 therapists
     14 therapy
      1 there
      1 thesis
      1 thess
      1 thessalien
      1 thessaliska
      1 thessalum
      1 thetaperioder
      5 thetavågor
      2 they
      1 th�ger
      1 thibetanus
      1 thick
      1 thiel
      2 this
      1 thjälparceller
      1 thjälparcellerna
      1 thjälparlymfocyter
      1 thoeris
      2 thom
     17 thomas
      2 thompson
      1 thomson
      1 thor
      1 thoracic
      1 thorax
      1 thoraxintensivvård
      1 thoraxkirurger
      3 thoraxkirurgi
      1 thoraxröntgen
      1 thoraxröntgenden
      1 thoraxskador
      1 those
      1 thought
      1 thpb
      1 thrane
      5 threading
      1 three
      1 threspons
      1 thriller
      1 throat
      1 thrombocytopenic
      1 thüringen
      1 thymol
      1 thymolum
      4 thymus
      1 thyreodit
      1 thyreoideastimulerande
      1 thyroarytenoidmuskeln
      5 thyroidea
      2 thyroideacancer
      1 thyroideae
      1 thyroideavävnad
      1 thyroidit
      1 ti�
      2 tia
      1 tiamin
      1 tiaminaserna
      1 tianbao
      1 tianjin
      7 tibast
      1 tibastbuskens
      1 tibastens
      1 tibastsläktet
      2 tibastväxter
      1 tibc
      1 tibern
      1 tiberön
      4 tibet
      2 tibetanska
      1 tibial
      1 tibialis
      1 tibialt
      1 tibiaperiostit
      1 tibiasyndrom
      1 tica
      1 tick
      1 ticka
      1 tickande
      1 tickborne
      4 tickor
     27 tics
      5 ticsen
    406 tid
      3 tidalvolym
      5 tidalvolymen
      2 tidbas
      2 tidbasen
      2 tidbasoscillatorn
      1 tidea
      1 tidelag
    180 tiden
      6 tidens
     41 tider
      3 tideräkning
      4 tiderna
      1 tidernas
      8 tiders
      1 tidevarv
     65 tidig
     89 tidiga
    371 tidigare
      6 tidigast
     15 tidigaste
      1 tidigmoderna
    174 tidigt
      1 tidlös
      4 tidlösa
      2 tidlösan
      1 tidlösasläktet
      1 tidlösasläktets
      3 tidlöseväxter
      1 tidlösor
      2 tidlösorna
      1 tidning
      5 tidningar
      1 tidningarna
      4 tidningen
      1 tidningsartiklar
      1 tidningsomslag
     20 tidpunkt
     10 tidpunkten
      6 tidpunkter
     24 tids
      1 tidsandar
      1 tidsaspekt
      1 tidsaspekten
      1 tidsåtgången
      2 tidsbegränsad
      2 tidsbesparande
      1 tidsbestämma
      1 tidsbokning
      1 tidscykler
      1 tidsdiagram
      1 tidsdomän
      1 tidsdomänens
      2 tidsenhet
      1 tidsfördröjande
      1 tidsförlopp
      1 tidsförloppet
      1 tidsfristen
      1 tidsgräns
      1 tidsinställd
      4 tidsintervall
      1 tidsintervaller
      1 tidsintervallet
      1 tidskänsliga
      4 tidskrävande
     10 tidskrift
     13 tidskriften
      4 tidskrifter
      1 tidskrifterna
     13 tidsperiod
      1 tidsperioden
      4 tidsperioder
      3 tidssamband
      1 tidsskalor
      1 tidsskillnad
      1 tidstypiska
      1 tidszon
      3 tidszoner
      1 tidtabeller
      1 tiemannspets
      1 tienlig
      1 tierno
      1 tiger
      1 tigermussling
      1 tigermusslingen
      1 tigersalamander
      1 tigersalamandern
      2 tight
      2 tighta
      1 tigrinus
      1 tikar
      1 tiken
      2 til
   8246 till
      1 tillaga
      2 tillagar
      1 tillagas
      5 tillagat
     12 tillägg
      1 tillägga
      2 tilläggas
      1 tilläggen
      1 tillägget
      1 tilläggs
      1 tilläggsavtal
      1 tilläggsbehandling
      1 tilläggsdiagnoser
      1 tilläggskost
      1 tilläggsskylt
      2 tilläggsspecialitet
      1 tilläggsspruta
      3 tilläggstavla
      1 tilläggstavlan
      1 tilläggstavlor
      1 tilläggstjänster
      2 tillägna
      1 tillägnad
      2 tillägnade
      4 tillagning
      3 tillagningen
      1 tillagningssätt
      1 tillagninguppvärmning
      8 tillämpa
      3 tillämpad
      2 tillämpade
      5 tillämpades
      1 tillämpande
      3 tillämpar
      1 tillämpare
     15 tillämpas
      1 tillämpat
      1 tillämpats
      2 tillämplig
      1 tillämpligt
     12 tillämpning
     19 tillämpningar
      2 tillämpningarna
      4 tillämpningen
      1 tillämpningsområden
      1 tillämpningsprocessen
      8 tillåta
      4 tillåtas
      1 tillåtelse
      1 tillåten
     33 tillåter
     23 tillåtet
      9 tillåtna
     12 tillåts
      3 tilläts
    123 tillbaka
      1 tillbakabildar
      4 tillbakabildas
      1 tillbakadragande
      2 tillbakadragandet
      2 tillbakadragen
      2 tillbakadragenhet
      1 tillbakadragningen
      5 tillbakagång
      1 tillbakahållande
      6 tillbaks
      2 tillbeds
      6 tillbehör
      1 tillblivelse
      1 tillbringa
      1 tillbringade
      5 tillbringar
      6 tillbud
      3 tilldelad
      1 tilldelade
      8 tilldelades
      1 tilldelar
      6 tilldelas
      1 tilldelning
      1 tilldrog
      1 tillerosa
      1 tillexo
     27 tillfälle
     29 tillfällen
      1 tillfällena
      8 tillfället
     37 tillfällig
     12 tillfälliga
      2 tillfällighet
      1 tillfälligheten
     41 tillfälligt
      2 tillfälligtvis
      1 tillfångatagen
      1 tillfångatagit
      1 tillflöde
      1 tillflödet
      1 tillflykt
      1 tillfoga
      1 tillfogar
      9 tillför
     15 tillföra
      5 tillföras
      3 tillförd
      1 tillförda
      6 tillförlitlig
      9 tillförlitliga
     10 tillförlitlighet
      1 tillförlitligheten
      5 tillförlitligt
     17 tillförs
      1 tillförsäkra
     21 tillförsel
      3 tillförseln
      3 tillfört
      2 tillförts
      3 tillfrågade
      1 tillfrågades
      2 tillfrån
      2 tillfreds
      2 tillfredsställa
     10 tillfredsställande
      8 tillfredsställelse
      1 tillfredsställer
      9 tillfriskna
      4 tillfrisknade
     11 tillfrisknande
      6 tillfrisknandet
      7 tillfrisknar
      4 tillfrisknat
      1 tillfriskningskvot
      8 tillgå
     51 tillgång
      5 tillgångar
      1 tillgångarna
     21 tillgången
     22 tillgänglig
     22 tillgängliga
      3 tillgänglighet
      6 tillgängligheten
     22 tillgängligt
      1 tillgick
      1 tillgivenhet
      1 tillgivenheten
      1 tillgjorda
      1 tillgodogjort
      6 tillgodogöra
      5 tillgodose
      2 tillgodosedda
      1 tillgodoser
      1 tillgripa
      2 tillgripas
      1 tillgriper
      1 tillgrips
      1 tillhåll
      5 tillhandahålla
      1 tillhandahållas
      8 tillhandahåller
      1 tillhandahålles
      2 tillhandahålls
    103 tillhör
      2 tillhöra
     23 tillhörande
      4 tillhörde
      1 tillhöriga
      1 tillhörighet
      2 tillhörigheter
      1 tillhörigt
      2 tillhört
      1 tillika
      1 tillintetgöra
      4 tillit
      1 tillitsfulla
      1 tillkalla
      1 tillkallade
      1 tillkallades
      1 tillkännagav
      1 tillkännagavs
      1 tillkännagifwande
      1 tillkännagivande
      1 tillkännagjorde
      5 tillkom
     10 tillkommer
      9 tillkommit
      1 tillkomna
      2 tillkomst
      1 tillkomsten
      1 tillnamn
      1 tillnyktringen
      1 tillo
      1 tillorsaka
      1 tillorycka
      1 tillpassa
      1 tillpassat
      1 tillpassning
      4 tillplattad
      1 tillplattade
      2 tillpressat
     31 tillräcklig
      8 tillräckliga
    120 tillräckligt
      1 tillräkneliga
      4 tillrätta
      2 tillredas
      1 tillreder
      1 tillredning
      3 tillreds
      1 tillretts
     82 tills
      1 tillsagd
    225 tillsammans
     19 tillsats
      1 tillsatsämnen
      4 tillsatsen
      8 tillsatser
      7 tillsatt
      3 tillsatta
     11 tillsätta
      1 tillsättas
      2 tillsatte
      5 tillsätter
      4 tillsattes
      3 tillsättning
      1 tillsättningen
      4 tillsatts
     14 tillsätts
      2 tillse
      1 tillskapas
      1 tillskillnad
      8 tillskott
      1 tillskrev
      3 tillskrevs
      1 tillskrivas
      1 tillskriver
      4 tillskrivits
      1 tillskrivna
      6 tillskrivs
      1 tillslutandet
      1 tillslutning
      1 tillslutningens
      1 tillsluts
      2 tillsmälta
    454 tillstånd
      1 tillståndbr
     12 tillstånden
    179 tillståndet
      2 tillstånds
      1 tillståndsavdelningen
      1 tillståndsdelen
      1 tillståndsgivande
      1 tillståndskrav
      1 tillståndsmaskin
      3 tillsvidare
     13 tillsyn
      2 tillsynen
      1 tillsynsavdelningen
      4 tillsynsmyndighet
      2 tillta
     12 tilltagande
      5 tilltal
      2 tilltala
      4 tilltalande
      1 tilltalas
      1 tilltalet
      2 tilltäppning
      1 tilltäppt
      2 tilltäppta
      5 tilltar
      1 tilltog
      4 tillträde
      1 tillträdesskydd
      4 tilltro
      1 tilltryckt
     10 tillvägagångssätt
      9 tillvägagångssättet
      4 tillvänjning
      1 tillvänjningen
      3 tillvara
      2 tillvarata
      1 tillvaratagande
      1 tillvaratar
      1 tillvaratas
      7 tillvaro
      9 tillvaron
      2 tillvarons
      6 tillväxa
     13 tillväxer
     54 tillväxt
      1 tillväxtcentrum
     27 tillväxten
      2 tillväxtfaktor
      7 tillväxtfaktorer
      1 tillväxtfaktorreceptor
      1 tillväxtfaktorreceptorn
      3 tillväxtfas
      1 tillväxtfasen
      1 tillväxtförlusten
      2 tillväxthämmande
      1 tillväxthastighet
      1 tillväxthastigheten
     35 tillväxthormon
      3 tillväxthormonbrist
      5 tillväxthormonet
      2 tillväxthormonets
      1 tillväxthormonfrisättande
      1 tillväxthormonnivåerna
      2 tillväxthormonproducerande
      1 tillväxtmönstret
      1 tillväxtperiod
      1 tillväxtreglering
      2 tillväxtspurt
      1 tillväxtstimulering
      1 tillväxttakt
      2 tillväxtzonerna
     37 tillverka
      9 tillverkad
     25 tillverkade
     16 tillverkades
      1 tillverkande
     22 tillverkar
     20 tillverkare
      7 tillverkaren
      1 tillverkarens
      8 tillverkarna
      1 tillverkarnas
     78 tillverkas
     12 tillverkat
     10 tillverkats
     47 tillverkning
     18 tillverkningen
      1 tillverkningsföretag
      1 tillverkningskedjan
      1 tillverkningsmetod
      1 tillverkningsprocessen
      1 tillverkningsprocessens
      1 tillverkningsprocesser
      1 tillverkningssed
      2 tim
      1 timberlake
      1 timbuktu
      6 time
      1 timediv
      1 timeoutmetoden
      2 timer
      3 times
      1 timglasfiguren
      1 timglasfigurer
      4 timglasformad
      1 timglasformade
      3 timing
      2 timjan
      1 timjankamfer
      1 timjanolja
    125 timmar
      1 timmar�
      1 timmarna
      8 timmars
     15 timme
      3 timmen
      2 timmes
      1 timor
      2 timori
      1 timotej
      1 timothy
      1 timrad
      1 tinar
      1 tinas
      1 tinats
     10 tinea
      1 tinells
      8 ting
      1 tingens
      1 tingest
      1 tingsrätt
      1 tingsrätten
      1 tinire
      1 tinktur
      1 tinktura
      1 tinkturer
      1 tinnar
      1 tinningbenets
      1 tinningen
      1 tinningloben
      1 tinninglober
      1 tinninglobernas
     63 tinnitus
      1 tinnitusartat
      1 tinnitusbesvären
      1 tinnitusdrabbade
      1 tinnitusen
      1 tinnitusklinikens
      1 tinnitusproblem
      1 tinnitussignalen
      1 tiny
     66 tio
      1 tiocyanat
      7 tionde
      2 tiondel
      1 tiondels
      2 tiopentalnatrium
      6 tiotal
      2 tiotals
      3 tiotusen
      1 tiotusendedel
      4 tiotusentals
      1 tiparol
      1 tipp
      2 tippar
      1 tippas
     10 tips
      1 tiptoe
      1 tirefond
      1 tirsa
      1 tirumalai
      2 tissue
      1 tistelfröolja
     11 titan
      1 titanbågar
      1 titandioxid
      1 titanet
      1 titanhakar
      1 titanvitt
      7 titel
      1 titelförsvararen
     19 titeln
      1 titelskydd
      1 titer
      1 titerstegring
      3 titlar
      1 titt
     11 titta
      1 tittade
     18 tittar
      1 tittarna
      1 tittarstorm
      2 tittat
      1 titthål
      4 titthålskirurgi
      1 titthålskirurgiskmetod
      2 titthålsoperation
      1 titthålsteknik
      1 tituleras
      1 tiva
      1 tjackballe
      1 tjackrace
      1 tjälen
      1 tjällossningstid
      1 tjäna
      1 tjänade
      4 tjänar
      3 tjänare
      1 tjänarna
      1 tjänat
      1 tjänlig
      1 tjänligt
      7 tjänst
      2 tjänstefel
      1 tjänstefolket
      5 tjänstehund
      2 tjänstehundar
      1 tjänstehundskort
      1 tjänsteman
      1 tjänstemän
      1 tjänsteorienterade
      1 tjänsteplikt
     12 tjänster
      1 tjänsteresor
      1 tjänsterna
      1 tjänstgjorde
      2 tjänstgör
      1 tjänstgöra
      4 tjänstgöring
      1 tjänstgöringarna
      5 tjära
      2 tjärfärgämnen
      1 tjäroljefraktion
      1 tjäror
      1 tjärpapp
      1 tjeckien
      1 tjeckiska
      1 tjeckiske
      2 tjeckoslovakien
      1 tjeckoslovakisk
      1 tjej
      2 tjejer
      1 tjenlig
      1 tjernobylolyckan
     18 tjock
     19 tjocka
      1 tjockända
     14 tjockare
      1 tjockhudad
      1 tjockhudade
      1 tjockisen
     10 tjocklek
      4 tjockleken
      1 tjockleksmätningar
     12 tjockt
      2 tjocktarm
     47 tjocktarmen
      2 tjocktarmens
      1 tjocktarmepitelet
      1 tjocktarmsbakterier
      4 tjocktarmscancer
      1 tjocktarmsinnehåll
      1 tjocktv
      1 tjockväggiga
     11 tjugo
      1 tjugoandra
      1 tjugofem
      1 tjugonde
      3 tjugotal
      1 tjugotals
      1 tjugotvå
      1 tjur
      1 tjurar
      1 tjurfäktning
      1 tjut
      1 tjuv
      1 tjuvar
      1 tjuvjakt
      1 tk
      2 tlc
      1 tlingiterna
      1 tlinglitstammarna
      1 tljuden
      1 tlll
      2 tlr
      3 tlv
      5 tlymfocyter
      5 tlymfocyterna
      2 tlymphotropic
      2 tm
      1 tma
      1 tmattp
      3 tmpsmx
      2 tnf
      1 tnfa
      1 tnfalfa
      2 tnm
      1 tnmklassifikation
      1 tnmstadieindelningssystemet
      1 tnmsystemet
     21 to
      1 toabesök
      8 toalett
      1 toalettartiklar
      5 toalettbesök
     11 toaletten
     10 toaletter
      1 toaletthandduk
      1 toaletthandduken
     10 toalettpapper
      6 toalettpapperet
      1 toalettpapperets
      1 toalettpappershållare
      1 toalettpapperstillverkarna
      1 toalettpappret
      1 toalettsaker
      1 toalettsits
      1 toalettsitsar
      4 toalettstolar
      3 toalettstolen
      1 toalettvanor
      1 töar
      1 töat
      3 tobacco
     51 tobak
      7 tobaken
      2 tobakens
      1 tobaksanvändning
      1 tobaksbehållare
      1 tobaksexportörer
      1 tobaksförbrukning
      1 tobaksförsäljare
      1 tobaksglöd
      1 tobaksindustrin
      1 tobakskalebasser
      1 tobakskonsumtionen
      1 tobaksodlingarna
      2 tobakspipor
      2 tobaksprodukter
      1 tobakspung
      1 tobakspungar
      2 tobaksransoner
      1 tobaksreklam
      1 tobaksrelaterade
      1 tobaksrevolutionen
      4 tobaksrök
      2 tobaksrökare
      1 tobaksröken
     12 tobaksrökning
      2 tobaksrökningen
      1 tobaksväxter
      1 tobias
      1 toe
      1 tof
      1 toffee
      2 toffelblomma
      1 tofflor
      1 tofs
      1 tofsar
      1 tofsskivlingar
      3 tofu
      2 tofus
     57 tog
      1 togo
     29 togs
      1 toivo
      1 töja
      3 töjas
      1 töjbara
      1 töjer
      2 töjning
      1 töjningen
      1 tokajer
      1 tokfursten
      1 tokig
      1 tokujiro
      2 tokyo
      1 tokyopolisen
      1 tokyos
      1 told
      1 tolerabilitet
      1 tolerance
      3 tolerans
      3 toleransen
      1 toleransnivån
      1 toleransökning
      3 toleransutveckling
      4 tolerera
      1 tolererar
      6 tolereras
      1 tolererat
      2 tolfte
     18 tolka
      2 tolkade
      2 tolkades
      1 tolkandet
     11 tolkar
      1 tolkaren
     20 tolkas
      1 tolkat
      4 tolkats
      1 tolkcentral
     20 tolkning
      7 tolkningar
      3 tolkningen
      1 tolkningsansvar
      1 tolkningsförslag
      1 tolkningsprocess
      1 tolkningstraditionen
      1 tolleen
      2 tolllike
      6 toluen
      1 toluensulfonamid
      1 toluol
     24 tolv
      1 tolvåriga
      1 tolvfinge
      1 tolvfingertarm
     28 tolvfingertarmen
      5 tolvfingertarmens
      1 tolvmånadersperiod
      2 tolvstegsprogram
      1 tolvstegsprogrammen
     13 tom
      4 tomas
      3 tomat
      1 tomaten
      2 tomater
      1 tomb
      1 tömbar
      2 tömd
      1 tömde
      4 tome
      2 tomentosum
      1 tomentosus
      1 tomhet
      2 tomma
     20 tömma
      6 tömmas
      7 tömmer
      1 tommy
     16 tömning
      2 tömningarna
      1 tömningen
      1 tomograf
      8 tomografi
      1 tomografin
      3 tomografisk
      2 tomografiska
      1 tomografitekniken
      1 tomogram
      2 tomography
      2 tomrum
     15 töms
      3 tomt
      1 tomtarm
      3 tomtarmen
      2 tomtebloss
      2 tömts
     27 ton
      1 �ton
      1 tonaccenter
     11 tonande
      1 tonår
     15 tonåren
      1 tonåriga
      9 tonåringar
      1 tonåringarna
      1 tonåringen
      2 tonårsflickor
      2 tonårsidol
      1 tonårsidoler
      2 tonaudiometri
      1 tondöv
      1 tonen
     10 toner
      1 tonerna
      1 toneurytmi
      1 toneurytmin
      2 tonfisk
      1 tongivare
      7 tonhöjd
      2 tonhöjden
      1 toning
      4 tonlägen
      9 tonlatens
      3 tonlatensen
      1 tonlatenstyper
      2 tonlatenstyperna
      5 tonlösa
      1 tonlöst
      2 tonometer
      1 tonometern
      1 tonometrar
      4 tonometri
      1 tonometriförfarandet
      1 tonsillerna
      4 tonsillit
     12 tonsilloliter
      1 tonskalan
      1 tonsurans
      1 tönt
      2 tonterapi
      1 töntig
      1 töntprylstämpel
      1 tontröskel
      3 tonus
      2 tonvikt
      1 tonvikten
      1 tony
      2 topf
      3 topfree
      4 topfreedom
      3 topiken
      1 topiska
     24 topless
      1 toplessaktioner
      2 toplessmodet
      2 toplesssolandet
      1 topografi
      2 topografiska
     12 topp
      3 toppar
      8 toppen
      1 toppidrottare
      1 toppigt
      1 toppkonsument
      1 topplöst
      3 toppmatad
      2 toppmatade
      1 toppmöten
      1 toppmötet
      1 topprider
      2 toppskikt
      5 toppställda
      1 topptio
      1 topsning
      1 tor
      1 torakala
      6 torakalt
      2 torakocentes
     12 torde
      1 törelsläktet
      3 törelväxter
      3 torg
      3 torgskräck
      6 torium
      1 toriumdioxid
      1 toriumreserver
      2 tork
     31 torka
      3 torkad
      6 torkade
      1 torkande
     14 torkar
      7 torkas
      2 torkat
      1 torkats
      2 torkel
      1 torklada
      1 torkladan
      1 torkladans
      2 torklina
      3 torkmedel
      1 torkmetod
      1 torkmetoder
      9 torkning
      1 torkprocess
      9 torkskåp
      1 torkskåpen
      1 torkstuga
      1 torktåliga
      7 torktumlare
      2 torktumlaren
      1 torktumling
      1 torkvinda
      1 törlarnas
      1 torminosus
      1 torn
      1 tornerspel
      1 tornet
      3 toronto
      1 torontos
      2 torparkex
      2 torpeder
      1 torquata
     23 torr
     24 torra
      1 torrare
      1 torrbastu
      3 torrbatterier
      1 torrdassen
      2 torrdestillation
      1 torrdiskning
      2 torrdräkt
      1 torrey
      1 torreyi
      1 torrfläcksjuka
      5 torrhet
      1 torrheten
      1 torrhetskänsla
      4 torrhosta
      2 torris
      1 torrisbehandling
      1 torrisen
      1 torrissnö
      1 torrlades
      1 torrlagda
      1 torrmjölk
      1 torröra
      2 torröta
      1 torrplåtenoch
      1 torrpreparat
      1 torrsättning
      2 torrschampo
      1 torrsubstanshalten
     12 torrt
      2 torrtiden
      2 torrvaror
      1 torrvikten
      1 torsdagskväll
      1 torseletter
      1 torshälla
      3 torsion
      1 torsite
      2 torsk
      4 torskmask
      1 torslanda
      1 torson
      1 torsson
     16 törst
      1 törstcentrum
      2 törsten
      1 törstig
      1 törstiga
      1 törstkänslorna
      4 torticollis
      1 tortyr
      1 tortyrredskap
      1 torulaspora
      1 torus
      1 torvbottnar
      1 toscana
      1 toshiba
      1 toshikazu
     36 total
     34 totala
      1 totalantalet
      1 totalbedövning
      1 totalbekämpningsmedel
      1 totalförbjudits
      1 totalförbud
      1 totalförsvarsplikt
      1 totalintravenös
      2 totalstopp
     29 totalt
      9 tourettes
      1 tourettsliknande
      1 �tournefortii
      1 tourniquet
      1 tourniquettest
      2 tourniquettestet
      1 tovar
      1 tovning
      1 towern
      1 townsite
      2 toxic
     11 toxicitet
      1 toxiciteten
      1 toxicitetsstudier
      4 toxicodendron
      1 toxicos
      1 toxikokinetik
      7 toxikologi
      1 toxikologin
      1 toxikologisk
      1 toxikologiska
      1 toxikon
     14 toxin
     16 toxiner
      4 toxinerna
     10 toxinet
      1 toxinets
      1 toxinhalterna
      1 toxinologi
      6 toxisk
     25 toxiska
      6 toxiskt
      1 toxitet
      1 toxocariasis
      1 toxoid
      1 toxoider
      5 toxoplasma
      1 toxoplasmaägg
      3 toxoplasmos
      2 toxorhynchites
      1 tp
      1 tpb
      1 tpn
      1 tpr
      1 tptid
      1 tr
     29 trä
      1 trabekulära
      4 träben
      1 träbenet
      2 träbit
      1 träbitar
      1 träbyggnad
      1 traces
      5 trachea
      1 trachealkanyl
      1 trachealkanylen
      2 tracheostoma
      1 tracheostomi
      6 trachomatis
      1 trachycarpus
      1 track
      1 tracy
      1 tracyi
      1 trad
      8 tråd
     44 träd
      2 träda
      1 trädansamlingar
     11 trådar
      1 trådarna
      1 trädart
      9 trädde
      1 träddes
      2 tråddragande
      1 trade
     12 tråden
      5 träden
      1 trädens
      2 träder
      8 trädet
      5 trädets
      1 trådformade
      2 trådformiga
      1 trädgård
     10 trädgårdar
      1 trädgården
      1 trädgårds
      1 trädgårdsformer
      1 trädgårdshandeln
      1 trädgårdsland
      7 trädgårdsväxt
      4 trädgårdsväxter
      1 trädgränsen
     24 tradition
      1 traditional
     23 traditionell
     38 traditionella
     34 traditionellt
      8 traditionen
      7 traditioner
      4 traditionerna
      1 trådlika
      1 trådliknande
      1 trådlös
      3 trådlösa
      1 trädnöts
      1 tradolan
      1 trädrot
      1 trådsmala
      1 trädstubbar
      1 trådtunna
      3 träet
      1 träets
      1 träff
     11 träffa
      2 träffades
     14 träffar
      3 träffas
      1 träffat
      1 träffens
      3 traffic
      5 trafik
      1 trafikanten
     12 trafikanterna
      4 trafikbuller
      1 trafikdödad
      1 trafikdödas
      4 trafiken
      2 trafikerade
      1 trafikerar
      1 trafikflygplan
      1 trafikmedicin
      1 trafikmiljön
      5 trafikolyckor
      1 trafikolyckorna
      1 trafiköverträdelser
      1 trafikpolis
      1 trafiksäkerhet
      2 trafiksignal
      1 trafiksignaler
      1 trafikslagen
      2 trafikverket
      1 tragusömhet
      1 trailer
      1 trails
      1 träimpregnering
      1 train
      2 training
      1 trakassera
      1 trakasserar
      1 trakasserier
      3 trakea
      1 trakealkanyl
      1 trakeostomi
      6 trakeotomi
      1 träklubba
      2 träkol
      2 trakom
      1 träkonstruktioner
      2 trakt
      2 trakten
      4 trakter
      2 trakterna
      1 traktorer
      1 tralala
      1 träls
      1 trälträlinna
      2 tramadol
      1 trampa
      1 trampat
      1 trampolinen
     25 träna
      2 tränad
      3 tränade
      1 tränande
     12 tränar
      2 tränas
      6 tränat
      3 tränats
      1 tranbär
      1 tranbärsjuice
      1 tranbärstillsats
      1 trance
      1 trancopal
      1 tranexamsyra
      8 trång
      6 trånga
     21 tränga
      2 trängande
      2 trångboddhet
      1 trångbott
      1 trängde
      1 trängdes
     18 tränger
      1 trängingsinkontinens
      1 trängning
      5 trängningsinkontinens
      2 trängre
      1 trängs
      4 trängsel
      2 trångt
      3 trängt
      1 trångvinkelglaukom
    103 träning
     14 träningen
      2 träningens
      4 träningsberoende
      4 träningsberoendet
      1 träningscyklar
      1 träningsdos
      1 träningsdosen
      1 träningsform
      1 träningsformen
      2 träningsformer
      1 träningsinducerad
      1 träningsinsats
      3 träningsintolerans
      1 träningsmetod
      1 träningsmetoder
      1 träningsnarkomani
      1 träningsområdet
      5 träningspass
      4 träningspasset
      1 träningspassets
      1 träningsperioden
      1 träningsperioder
      5 träningsprogram
      1 träningsreglering
      1 träningsskola
      1 träningssystem
      2 träningsvärk
     12 trans
      5 transactional
      2 transaktioner
      5 transaktionsanalys
      7 transaktionsanalysen
      1 transaktionsanalysens
      6 transaktionsanalytiker
      4 transaktionsanalytikern
      1 transaktionsanalytiska
      1 transaktionsanlysen
      2 transaminaser
      1 transaminaserna
      1 transanal
      1 transartat
      1 transavia
      2 transcendenta
      1 transcendental
      1 transcendentalists
      3 transdermala
      1 transdermalt
      1 transducer
      1 transe
      2 transen
      1 transendotelisk
      1 transesofageal
      1 transfer
      1 transferasbrist
      4 transferrin
      1 transferrinbestämning
      1 transferrinbundet
      1 transferrinet
      1 transferrinkomplex
      1 transferrinmättnad
      1 transferrinreceptorer
      1 transferrinvärde
      5 transfetter
      5 transfettsyror
      1 transfixation
      2 transformation
      1 transformator
      1 transformeringen
      2 transforming
      5 transfusion
      1 transfusionen
      5 transfusioner
      1 transfusionsreaktioner
      1 transfusionssmitta
      1 transglutaminaser
      1 transglutaminaset
      1 transglutminas
      1 transient
      1 transientskyddad
      1 transire
      1 transisomer
      1 transistorer
      1 transistorerade
      1 transithamnarna
      1 transitions
      2 transitorisk
      2 transkortikal
      1 transkriberas
      1 transkriberat
      1 transkript
      2 transkriptas
      1 transkription
      6 transkriptionen
      1 transkriptionsfaktorer
      3 transkutan
      1 translationell
      1 translationen
      1 transliknande
      3 translokation
      1 translokationer
      1 translokeringssteget
      1 transluminal
      1 transluminell
      1 transmembrana
      1 transmembranreceptor
      1 transmissionsvägen
      1 transmittorsubstansen
      3 transmittorsubstanser
      1 transmural
      2 transmutation
      1 transmuteras
      1 transparensforum
      5 transparent
      1 transparenta
      1 transpeptidasenzym
      1 transpeptidasenzymerna
      1 transpeptidasenzymet
      1 transpeptideringnsreaktionen
      1 transpeptideringsreaktionen
      1 transperson
      1 transpersonell
      1 transpersonella
      1 transpersoner
      1 transpiration
      4 transplantat
      1 transplantaten
      1 transplantatet
     18 transplantation
      6 transplantationer
      1 transplantationerna
      1 transplantationsförsök
      1 transplantationskirurgin
      1 transplantatmotvärdsjukdom
      3 transplantera
     14 transplanterade
      3 transplanteras
      1 transpolyisopren
     14 transport
      1 transportalternativ
      4 transporten
      1 transportepitel
      3 transporter
     18 transportera
     16 transporterar
     42 transporteras
      1 transporterna
      1 transportföretaget
      1 transportförmåga
      1 transportglobulin
      2 transportkanaler
      2 transportmedel
      1 transportmöjligheterna
      1 transportör
      1 transportören
      4 transportprotein
      3 transportproteiner
      4 transportsystem
      1 transposoner
      1 transpotera
      3 transsexualism
      1 transsexuell
      4 transsexuella
      1 transsfenoidal
      1 transställning
      1 transsudat
      2 transthyretin
      7 transtillstånd
      1 transtorakal
      1 transtorakalt
      1 transuran
      1 transuranen
      1 transuraner
      1 transversal
      1 transversalplanet
      1 transversell
      2 transversus
      1 trap
      1 träplankor
      1 trappades
      3 trappor
      1 trappsteg
      2 trär
      1 träracketar
      1 träram
      1 träramar
      1 trare
      1 trärör
      2 träs
      4 trasa
      1 trasan
      1 trasig
      1 trasiga
      1 träslag
      1 träslaget
      1 träsnitt
      3 trasor
      1 träspatel
      1 träspjut
      4 träsprit
      1 trassla
      1 trastar
      1 trästicka
      1 tratt
      1 trätt
      1 trattar
      7 trattbröst
      1 trattbröstoperationer
      1 trattbröstpatienter
      1 trattformat
      1 trattlika
      1 trauer
     44 trauma
      1 traumaband
      1 traumabehandlingen
      1 traumaenheterna
      1 traumafokuserad
      1 traumahundar
      9 trauman
      1 traumarelaterade
      1 traumas
      1 traumata
      1 traumateam
      1 traumatic
      1 traumaticin
      1 traumatiserade
      7 traumatisk
     12 traumatiska
      1 traumatiskt
      5 traumatologi
      5 traumatologin
      3 traumdeutung
      1 trautmann
      1 träväggarna
      2 travail
      1 travell
      2 traverslyftar
    425 tre
      1 trea
      3 treårig
      2 treåriga
      2 treårigt
      1 treåring
      1 treårsåldern
      1 treårsperiod
      1 treating
      2 treatise
      5 treatment
      1 treblinka
      1 tredagars
      1 tredagarsbehandling
      1 tredagarskur
      3 tredelad
      1 tredelade
      1 tredelning
      1 tredimensionell
      7 tredimensionella
      3 tredimensionellt
     81 tredje
     22 tredjedel
      5 tredjedelar
      4 tredjedelen
      1 tredjedels
      1 tredrogsvarianten
      1 treenigheten
      1 trefaldig
      1 trefin
      1 treflikigt
      2 trefyra
      1 tregradig
      2 trehundra
      4 trekantig
      1 trekantiga
      1 treks
      2 trematoda
     13 tremens
      3 tremolit
      1 tremolitasbest
      1 tremolsianus
      4 tremor
      1 trenaunay
      1 trend
      3 trenden
      4 trender
      1 treo
      3 trepan
      1 trepanatio
      8 trepanation
      1 trepanationen
      1 trepanerad
      3 trepanerade
      2 trepanering
     16 treponema
      1 treponemaantikroppstest
      2 treponemal
      1 treponemaorsakade
      1 treponematest
      1 treponematester
      1 treponematoses
      2 treprocentig
      2 treschow
      1 treshold
      1 tresiffriga
      2 trettio
      1 trettioårsåldern
      3 trettiotal
      1 trettiotre
      4 tretton
      3 trevärd
      1 trevärda
      1 trevärt
      1 treves
      1 trevlig
      1 trevligare
      2 trevligt
      2 trh
      7 tri
      1 tria
      1 triacylglycerider
      2 triaden
      5 triage
      1 trial
      1 trials
      2 triangel
      1 triangelformad
      2 triangelformade
      1 triangulära
      1 triatominae
      1 triazin
      1 triazinring
      1 triazintriamin
      1 tribromresorcinol
      1 tribus
      1 tributyltenn
      2 tributyltennhydrid
      1 trich
      1 trichina
      7 trichinella
      1 tricho
      1 trichobilharzia
      3 tricholoma
      1 tricholomataceae
     12 trichomonas
      4 trichophyton
      1 trichorgaboutskinpickinghtml
      1 trichosanthes
      2 trichotillomani
      3 tricyklika
      2 tricyklisk
      8 tricykliska
      1 trier
      1 trierucateglyceroltrioleat
      2 trifokala
      1 trigeminus
      1 trigeminusnerven
      5 trigeminusneuralgi
      4 trigga
      3 triggade
      1 triggande
      7 triggar
      8 triggas
      1 triggbrus
      1 trigger
      1 triggern
      4 triggerpunkter
      1 triggsignal
      1 triglycerid
      5 triglycerider
      1 triglycerol
      3 trihalometan
      1 trijodmetan
      8 trijodtyronin
      1 trikå
      1 trikala
      1 trikinellainfektion
      1 trikinen
      6 trikiner
      1 trikininfektion
      1 trikinlarver
      9 trikinos
      1 triklina
      1 triklorättiksyra
      1 triklorbis
      1 trikloreten
      2 trikloretylen
      1 triklorhydroxidifenyleter
      3 triklormetan
     27 triklosan
      1 triklosans
      5 triklosantandkräm
      1 trikomonas
      1 trikomonaskolpit
      1 trikotillofagi
      9 trikotillomani
      2 trikuspidalklaffen
      1 trilla
      1 trillades
      2 trillingar
      1 trillingnerven
      1 trillingnervens
      1 trilux
      1 trimer
      2 trimestern
      7 trimetoprim
      1 trimetoprimsulfametoxasol
      3 trimetoprimsulfametoxazol
      1 trimetylamin
      1 trimetylaminuri
      1 trimetylentrinitramin
      2 trimix
      1 trimmat
      1 trimning
      1 trinitroresorcin
      1 trinukleotiden
      1 triol
      1 trioleate
      1 tripp
      2 trippeldiagnostik
      1 trippelkombination
      1 trippelnegativa
      1 trippelvaccin
      1 trips
      1 tripsis
     15 trisomi
      4 trisomier
      1 trisomierna
      1 trisomiformer
      1 trisomin
      1 tritagonist
      1 tritagonisten
      1 triumfer
      1 trivalenta
      1 trivalnamn
      1 trivas
      1 trivia
      7 trivialnamn
      2 trivialnamnet
     32 trivs
      2 trivseln
      1 trna
      1 trnamolekyler
      1 trnamolekylerna
     28 tro
      1 troa
      1 troakar
      1 trochanterbälte
      1 trockenbeerenauslese
      1 troctomorpha
      1 tröd
      1 trodd
     34 trodde
      5 troddes
      1 troende
      1 troeng
      1 troféer
      1 trofinivå
      1 trofoblaster
      1 trofoblasterna
      1 trofozoit
      2 trofozoiten
      1 trög
      1 trögare
      6 trögflytande
      1 tröghet
      1 trögt
      3 trohet
      1 troheten
      1 troilius
      1 troja
      4 tröja
      1 tröjan
      1 tröjor
      1 tröjorna
      3 trolig
      2 troliga
      1 troligare
      2 troligast
      1 troligaste
     68 troligen
     15 troligt
     12 troligtvis
      2 trollbär
      1 trolldeg
      1 trolldom
      1 trolldruva
      1 trolldryck
      1 trollen
      1 trolleritrick
      1 trolli
      2 trollkarl
      1 trollkarlar
      1 trollkonst
      2 trollkunniga
      1 trollpåsar
      2 trolltrumman
      1 trollved
      2 trolovade
      1 trolovningen
      1 tromb
      1 trombektomi
     11 trombin
      1 trombocytens
     19 trombocyter
      5 trombocyterna
      3 trombocyternas
      1 trombocyters
      2 trombocytopen
     11 trombocytopeni
      1 trombocytopenisk
      1 trombocytplugg
      1 tromboelastografi
      2 tromboembolism
      2 trombofili
      6 tromboflebit
      1 tromboflebiten
     14 trombolys
      1 trombolytiskt
     11 trombos
      1 trombosen
      4 tromboser
      1 tromboserna
      1 trombosrubbning
      1 trombossjukdom
      2 trombotisk
      1 trombotiska
      3 trombyl
      1 trompe
      2 tromsöloka
     13 tron
      1 trondheim
      1 tropanalkaloid
      1 tropanalkaloiderna
      1 trophe
      1 tropical
      1 tropicalandinus
      2 tropikerna
      1 tropikfärg
      5 tropisk
     26 tropiska
      2 troponin
      1 troponiner
      1 troposmi
     83 tror
     68 tros
      2 trosa
      1 trosan
      1 tröskel
      3 tröskelvärde
      1 tröskelvärdesmodell
      2 trösklar
      1 trösklarna
      1 trosorna
     10 trosskydd
      1 trosskyddet
      2 tröst
      1 tröstande
      1 tröstlös
      1 trosuppfattning
    200 trots
      1 trotsåldern
      1 trotsande
      2 trotsiga
      2 trotsigt
     11 trotssyndrom
      7 trott
     11 trött
      3 trötta
      1 tröttande
      1 tröttare
      1 tröttcellulit
     96 trötthet
      4 tröttheten
      1 trötthetskänsla
      1 trötthetskänslor
      1 trötthetssymtom
      2 trötthetssyndrom
      1 trottoarkanter
      1 trousseaus
      1 trovärdighet
      1 trovärdigt
      2 troy
      7 trt
      3 trubbiga
      2 trubbigt
      1 trubbkantig
      1 truck
      1 trumbo
      1 trumbull
      7 trumhinnan
      1 trumhinneperforation
      2 trumma
      6 trumman
      1 trummandet
      1 trummor
      1 trumpeten
      1 trumpinnefingrar
      2 truncus
      1 trupp
      3 trupperna
      1 truppförflyttningar
      1 trupps
      1 truppslagsfärg
      1 trust
      1 truth
    111 tryck
     25 trycka
      1 tryckaccenter
      1 tryckande
      1 tryckarna
      2 tryckas
      2 tryckbandage
      1 tryckblåsan
     21 trycker
      1 tryckeri
     74 trycket
      1 tryckfallsjuka
     14 tryckfallssjuka
      1 tryckförändring
      1 tryckförändringar
      2 tryckförändringen
      4 tryckförband
      1 tryckgradient
      1 tryckgradienten
      2 tryckimpregnera
      1 tryckimpregnering
      1 tryckkabin
      1 tryckkammarbehandling
     10 tryckkammare
      3 tryckkammaren
      1 tryckkammarverksamheten
      1 tryckkänsla
      1 tryckkänsliga
      1 tryckknapp
      1 tryckknappar
      1 tryckkokare
      1 tryckkokning
      1 tryckömhet
      1 tryckpåverkan
      1 tryckreducering
      9 trycks
      3 trycksänkande
      1 trycksänkning
      1 trycksänkningar
      1 trycksänkningen
      1 trycksänkningssituationer
      1 trycksår
      1 trycksätta
      1 trycksättas
      1 trycksensorer
      1 tryckskillnad
      3 tryckskillnaden
      1 tryckskillnader
      1 tryckskillnadsskador
      1 tryckstegringen
      3 tryckstyrd
      8 tryckt
      2 tryckta
      2 tryckte
      1 trycktes
      1 trycktyngd
      1 tryckunderstödd
      1 tryckvågor
      1 tryckvågorna
      1 tryckvågsbehandling
      9 trygg
      3 trygga
      6 trygghet
      1 tryggheten
      1 trygghetsbehov
      1 trygghetsboende
      1 trygghetssökande
      3 tryggt
      1 trypanon
     14 trypanosoma
      3 trypanosomer
      2 trypanosomiasis
      2 trypsin
      1 trypsininhibitorer
      2 trypsinogen
      1 tryptamin
      1 tryptas
      1 tryptizol
      4 tryptofan
      1 ts
      1 tsaren
      1 tsarryssland
      1 tscore
      1 tsesnabbtester
      1 tsetse
      6 tsetseflugan
      3 tsetseflugor
      1 tsetseflugorna
     21 tsh
      1 tshirtar
      1 tshirtbh
      1 tshirts
      1 tshvärden
      1 tsp
      1 tsprit
      2 tsqaltubo
      1 tsqaltubodistriktet
      6 tss
      1 tsstoxin
      1 tsta
      1 tstac
      1 tstae
      1 tstao
      1 tstap
      1 tsvet
      1 tswana
      1 tsyndrom
      1 ttae
      2 tte
      1 ttg
      1 ttillgå
      2 ttm
      1 ttp
      6 tub
      1 tubdykning
      4 tuben
      2 tubens
      3 tuber
     28 tuberculosis
      1 tuberkelbacillen
      4 tuberkelbaciller
      1 tuberkelbacillers
      7 tuberkelbakterien
      1 tuberkelbakterier
      1 tuberkelbakterierna
      1 tuberkler
      1 tuberklerna
      1 tuberkulin
      1 tuberkulinprov
      3 tuberkulintest
      1 tuberkuloid
      1 tuberkuloida
    172 tuberkulos
      2 tuberkulosbakterier
      1 tuberkulosbehandling
      1 tuberkulosbehandlingen
      2 tuberkulosen
      1 tuberkulosepidemi
      2 tuberkulosfall
      4 tuberkulosfallen
      1 tuberkulosförekomsten
      1 tuberkulosformerna
      1 tuberkuloskontrollprogram
      1 tuberkuloskontrollstrategi
      6 tuberkulosmeningit
      1 tuberkulosodling
      1 tuberkulosoffer
      2 tuberkulospatienter
      1 tuberkulospatienternas
      1 tuberkulosrisk
      2 tuberkulosrisken
      1 tuberkulossjuka
      2 tuberkulossjukdom
      1 tuberkulossjukes
      6 tuberkulossmitta
      1 tuberkulossmittade
      1 tuberkulossmittor
      1 tuberkulossusceptibilitet
      2 tuberkulossymtom
      1 tuberkulosundersökning
      3 tuberkulosvaccin
      1 tuberkulosvaccinet
      1 tuberkulosvarianter
      2 tuberna
      1 tuberös
      1 tubulär
      1 tubulära
      1 tubule
      2 tubuli
      1 tubus
      1 tudelade
      3 tugg
      3 tugga
      1 tuggade
      2 tuggapparaten
      6 tuggar
      3 tuggas
      1 tuggmuskler
      2 tuggmusklerna
      2 tuggning
      2 tuggningen
      1 tuggsvårigheter
      1 tuggsystemet
      1 tuggtobak
      1 tuggummi
      1 tukhtensis
      1 tuktas
      1 tuktigt
      1 tulare
      2 tularemi
      4 tularensis
      1 tulipa
      1 tullen
      1 tulo
      1 tulpansläktet
      1 tum
      1 tumefaciens
      1 tummas
      2 tumme
      1 tummelisa
      6 tummen
      2 tummens
      1 tummoffer
      1 tumnagel
      3 tumor
     63 tumör
      1 tumörartad
      1 tumörbehandling
      1 tumörbildning
      4 tumörcell
      1 tumörcellen
     18 tumörceller
      5 tumörcellerna
      1 tumörcellsomvandling
      1 tumördoser
     88 tumören
     11 tumörens
    134 tumörer
     12 tumörerna
      1 tumörernas
      1 tumörers
      1 tumörfamilj
      1 tumörformen
      1 tumörframkallande
      1 tumörhålan
      1 tumörinvasion
      1 tumörkirurgi
      1 tumörklassifikation
      1 tumörlika
      1 tumörliknande
      4 tumörmarkör
      1 tumörmarkören
      3 tumörmarkörer
      1 tumörmassa
      2 tumörmassan
      1 tumörmisstanke
      1 tumörnekrosfaktor
      1 tumörnekrosfaktoralfa
      1 tumörnekrosfaktorer
      4 tumörområdet
      2 tumörs
      6 tumörsjukdom
      9 tumörsjukdomar
      1 tumörsjukdomen
      1 tumörstället
      1 tumörstorleken
      1 tumörsuppressiva
      1 tumörsuppressogen
      1 tumörsuppressorgen
      4 tumörsuppressorgener
      1 tumörsuppressorgenerna
      3 tumörtillväxt
      1 tumörtillväxten
      2 tumörtyp
      3 tumörtypen
      3 tumörtyper
      1 tumörtypers
      1 tumörutredningar
      1 tumörvarianter
      2 tumörvävnad
      1 tumörväxt
      1 tumörväxten
      3 tumregel
      1 tumregeln
      1 tumroten
      1 tumsidan
      7 tung
     32 tunga
     51 tungan
     13 tungans
      1 tungbenen
      1 tungbenet
      1 tungbett
      3 tungmetall
      8 tungmetaller
      1 tungmetallerna
      1 tungmetallförgiftning
      2 tungmusklerna
      1 tungor
      1 tungpiercing
      1 tungpiercingen
      1 tungrotenbr
      1 tungsinthet
      1 tungskrapa
      1 tungskrapan
      2 tungspat
      1 tungspetsenbr
      4 tungt
      1 tungviktsboxaren
      2 tunica
      1 tunika
      1 tunmören
     30 tunn
     23 tunna
      1 tunnar
     14 tunnare
      1 tunnas
      1 tunnaste
      4 tunnel
      1 tunnelbana
      3 tunneln
      3 tunnelseende
      1 tunnflytande
      2 tunnhåriga
      1 tunnskiktsdatortomografi
      1 tunnskiktskromatografi
      1 tunnslipad
      4 tunntarm
      1 tunntarmarna
     49 tunntarmen
     12 tunntarmens
      1 tunntarmsbiopsin
      2 tunntarmscancer
      1 tunntarmscellerna
      1 tunntarmssjukdom
      1 tunntarmsslynga
      1 tunntarmssvikt
      1 tunntarmstumörer
      1 tunnväggiga
     12 tunt
      2 tuppar
      1 tuppaskinn
      1 tuppkamsextrakt
      2 tupplur
      3 tupplurar
      2 tupplurarna
    142 tur
      2 turbin
      1 turbiner
      1 turbuhaler
      1 turbulenta
      2 turcica
      1 turer
      2 turism
      1 turistattraktion
      2 turistdiarré
      3 turister
      1 turistmål
      1 turistorten
      2 turkar
     13 turkiet
      1 turkiets
      1 turkiska
      1 turkos
      1 turksadeln
      1 turner
      3 turners
      1 tuschfärgning
     21 tusen
      1 tusenårig
      1 tusende
      2 tusendels
      1 tusenmoder
      1 tusental
     15 tusentals
      1 tuskaft
      1 tuskaftsvävd
      3 tuskegee
      1 tuskegeestudien
      4 tussilago
      2 tussilagon
      2 tussilagons
      1 tussipekt
      1 tussis
      1 tuta
      1 tutti
      1 tuukka
      1 tuulse
      1 tuva
      1 tuvad
      1 tuvade
     12 tv
    755 två
      4 tvåäggstvillingar
      4 tvåårig
      1 tvååriga
      1 tvåårsperiod
      1 tvåbasiga
      1 tvåbenta
      2 tvåbetygsnivån
      5 tvåbyggare
      1 tvådelad
      3 tvådimensionell
      2 tvådimensionella
      1 tvåfärgade
      1 tvåg
      4 tvågen
      2 tvågens
      4 tvagning
      3 tvågor
      1 tvågorna
      1 tvåhjärtbladiga
      1 tvåhjuligt
      2 tvåhundra
      1 tvåhundratalet
      1 tvåkärniga
      3 tvåkönade
     47 tvål
      1 tvåla
      1 tvålanvändning
      2 tvålar
      1 tvålbolags
     10 tvålen
      1 tvålframställning
      1 tvålliknande
      1 tvållösningar
      1 tvålopera
      1 tvålrester
      1 tvålsten
      2 tvåltillverkaren
      2 tvålvatten
      8 tvång
      3 tvånget
      6 tvångsbeteenden
      3 tvångsbeteendet
      1 tvångsförvaltning
      1 tvångshandling
      5 tvångshandlingar
      1 tvångshandlingarna
      2 tvångshandlingen
      1 tvångsimpulsiva
      1 tvångsintagna
      1 tvångsintagning
      6 tvångsmässig
      4 tvångsmässiga
      9 tvångsmässigt
      1 tvångsmedicinering
      1 tvångsrörelser
      2 tvångssteriliserades
      8 tvångssterilisering
      6 tvångssteriliseringar
      1 tvångssteriliseringarna
      1 tvångssteriliseringen
      1 tvångssymptomen
     37 tvångssyndrom
      7 tvångstankar
      4 tvångstankarna
      2 tvångstanke
      5 tvångstanken
     10 tvångsvård
      1 tvångsvis
      1 tvåpartssamtal
      1 tvåportsnätverk
      2 tvapparater
      1 tvapparaterna
      1 tvåprocent
      2 tvär
      1 tvära
      1 tväravbitare
      2 tvärbundna
      1 tvärdet
      1 tvärdrag
      3 tvären
      3 tvärgående
      1 tvärkulturella
      1 tvärled
      1 tvärrandningar
      1 tvärs
      1 tvärsnittsbild
      2 tvärsnittsstudie
      1 tvärsnittsstudier
      1 tvärsnittstudie
      1 tvärsnittyta
      2 tvärstrimmig
      2 tvärstrimmiga
      9 tvärt
      3 tvärtemot
     14 tvärtom
      1 tvårummig
      5 tvärvetenskaplig
      5 tvärvetenskapligt
      1 tvåstegsmetod
      1 tvåstegsprocess
      2 tvåtre
     34 tvätt
     26 tvätta
      2 tvättad
      1 tvättade
      2 tvättades
      1 tvättande
      9 tvättar
      1 tvättarbetet
      1 tvättarfamiljen
      1 tvättarfamiljs
     19 tvättas
      1 tvättat
      2 tvättats
      1 tvättbara
      1 tvättbart
      1 tvättbehandling
      1 tvättbiträde
      1 tvättbjörn
      2 tvättboll
      3 tvättbollar
      2 tvättbräda
      3 tvättbrädan
      1 tvätteffektivitetsklass
     11 tvätten
      1 tvätteri
      3 tvätterimuseum
      1 tvätterska
      1 tvättförkläden
      2 tvättgodset
      1 tvätthoar
      1 tvättid
      1 tvättkorgen
      1 tvättmadam
     19 tvättmaskin
      8 tvättmaskinen
      3 tvättmaskiner
      1 tvättmaskinerna
     13 tvättmedel
      1 tvättmedelsfack
      1 tvättmedlet
      1 tvättmetod
      1 tvättmetoder
      2 tvättmöjligheter
      5 tvättning
      1 tvättningrensning
      1 tvättpåsar
      2 tvättpelare
      1 tvättprogrammet
      1 tvättritualer
      3 tvättstuga
      1 tvättstugan
      3 tvättstugor
      2 tvättsvamp
      1 tvättsvampar
      1 tvättsymboler
      1 tvättverksamheten
      1 tvåtusen
      1 tvåvägs
      1 tvåvägsprocesser
      1 tvåvåningsbastun
      3 tvåvärd
      1 tvåvärda
      1 tvåvärt
      1 tvåveckorslinser
      1 tvåveckorsperiod
      1 tvåvingade
      2 tvåvingar
      1 tvbildrör
      2 tvbolaget
      1 tveeggad
      1 tvekade
      1 tvekan
      4 tveksam
      2 tveksamhet
      2 tveksamma
      4 tveksamt
      1 tvetydig
      2 tvetydiga
      1 tvhändelsen
      1 tvilling
      9 tvillingar
      1 tvillingarna
      1 tvillingbrodern
      2 tvillingbror
      1 tvillingen
      1 tvillinggraviditeter
      1 tvillingskaran
      5 tvillingstudier
      1 tvillingstudiers
      3 tvinga
      1 tvingad
      1 tvingade
      3 tvingades
      2 tvingande
      8 tvingar
     11 tvingas
      3 tvingats
      1 tvinnad
      2 tvinnade
      1 tvinnknut
      1 tvistar
      2 tvivelaktig
      1 tvivelaktiga
      1 tvivelaktigt
      1 tvivla
      1 tvivlar
      1 tvkanalen
      1 tvmärket
      1 tvprogram
      1 tvprogramledaren
      3 tvprogrammet
      1 tvradio
      2 tvserie
      3 tvserien
      2 tvserier
      3 tvskärm
      1 tvskärmen
      4 tvspel
      1 tvtittande
      6 tvungen
      3 tvungna
      1 twätt
      1 tweaking
      1 tweed
      2 twigg
      1 twin
      1 twinrix
      1 twoway
      1 tx
      4 ty
      6 tycka
      5 tyckas
      2 tycke
     25 tycker
     49 tycks
      7 tyckte
      1 tycktes
      1 tyd
     24 tyda
      1 tydde
     53 tyder
     30 tydlig
     22 tydliga
      9 tydligare
      7 tydligast
      1 tydligaste
      2 tydligen
      1 tydliggör
     48 tydligt
     12 tyfoidfeber
      7 tyfus
      1 tyfuspatienter
      1 tyfussjukdom
      1 tyfussjukdomar
     16 tyg
      1 tygband
      1 tygbindan
      6 tygbindor
      1 tygbit
      1 tygbörs
      5 tyger
      4 tyget
      1 tygfodral
      1 tyglager
      1 tyglande
      1 tyglar
      1 tygliknande
      1 tygremsa
      1 tygremsan
      1 tygstycke
      1 tygstycken
      1 tygtrosskydden
      1 tyler
      1 tyllbroderier
      1 tymidin
     10 tymol
      1 tymolförening
      1 tymolnatrium
      1 tympani
      1 tymushormoner
      2 tynade
      1 tyne
      1 tyngas
      1 tyngd
      1 tyngdkänslor
      1 tyngdlyftare
      3 tyngdpunkten
     12 tyngre
      1 tyngsta
    423 typ
      1 typart
      1 typdiabetes
      3 type
     63 typen
    290 typer
     22 typerna
      1 typfall
      1 typherix
      1 typhii
      1 typhim
      1 typhoidea
     15 typisk
     59 typiska
     54 typiskt
      1 typologi
      1 typsnitt
      1 tyr
      1 tyramin
      1 tyreglobulinet
      7 tyreoglobulin
      5 tyreoglobulinet
      1 tyreoidahormoner
      1 tyreoideahormon
      6 tyreoideahormoner
      2 tyreoideahormonerna
      1 tyreoideastimulerande
      1 tyreoidit
      2 tyreoperoxidas
      1 tyreoperoxidasen
      2 tyreotoxikos
      2 tyreotoxisk
      1 tyreotropinreceptorer
      1 tyreotropinreceptorerna
      1 tyrodeahormonerna
      2 tyroidea
      2 tyroideahormoner
      7 tyrosin
      3 tyrosinas
      1 tyrosine
      1 tyrosinet
      1 tyrosinkinas
      1 tyrosinkinase
      1 tyrosinkinastyp
      1 tyrotoxisk
      9 tyroxin
      2 tyroxinbindande
      1 tyroxinvärdet
      8 tysk
     34 tyska
      2 tyskamerikanska
      2 tyskan
      6 tyskans
      2 tyskarna
      1 tyskarnas
      1 tyskblodiga
     18 tyske
      4 tysken
     55 tyskland
      1 tysklands
      1 tysklönn
      3 tyskt
      1 tyson
      4 tyst
      5 tysta
      2 tystare
      1 tystlåtet
      2 tystnad
      7 tyvärr
      1 tzay
      1 tzeltalmayaner
     25 u
      1 ud
      1 udda
      1 uddbladet
      1 udden
      1 uddevalla
      1 uddspets
      1 uddspetsga
      1 udpavgår
      1 udpglukopyrufosforylas
      1 udpglukos
      1 udpglukosmolekylen
      1 udpglukosmolekyler
      1 ueshiba
      2 uet
      1 ufficiali
      2 uformad
      1 uformat
     15 uganda
      1 ugandas
      1 ugandisk
      1 ugandiska
      1 ugarte
      1 uggla
      1 uggleutgåvan
      1 ugglor
      1 ugn
      1 ugnen
      1 ugnsluckor
      1 ugnsrengöring
      1 ugnssteker
     10 uicc
      1 uiccs
      1 uitto
      1 uk
      1 ukärnorna
      6 ukraina
      1 ukrainetz
      6 uländer
      1 ulceration
      7 ulcerös
      7 ulcus
      1 ulf
      1 ull
      4 ulla
      1 ullånger
      1 ullen
      1 ullens
      1 ulleråkers
      1 ullig
      1 ullman
      1 ullöss
      1 ulm
      1 ulnaris
      1 ulnartunnelsyndrom
      1 ulrichii
      1 ulrik
      2 ulrika
      1 ultaljud
      1 ultimat
      1 ultimata
      1 ultra
      1 ultrabasiska
     32 ultraljud
      1 ultraljudsapparater
      1 ultraljudsbaserad
      2 ultraljudsbilder
      1 ultraljudscaler
      2 ultraljudsgivare
      3 ultraljudsgivaren
      3 ultraljudsteknik
      1 ultraljudstekniken
     14 ultraljudsundersökning
      3 ultraljudsundersökningar
      7 ultraviolett
      4 ultravioletta
      2 ulv
      1 ulvar
      1 ulvatand
      1 umami
      1 umas
      1 umbelliferon
     21 umeå
      1 umeälvens
      1 umeåregionen
     16 umgänge
      1 umgängesgrupp
      1 umgängesregler
      2 umgänget
      2 umgås
      1 umgicks
      1 umhlanga
      2 unaids
      1 �unconscious
      2 und
     31 undan
      1 undanhållas
      1 undanhålls
      1 undanråds
      2 undanröja
      1 undanröjs
      1 undanskymda
     47 undantag
      1 undantagen
      9 undantaget
      3 undantagna
      1 undantagsbestämelser
      3 undantagsfall
      1 undantagsregler
      1 undantagsvälde
      6 undantagsvis
      1 undantryckta
   2132 under
      1 underaktivitet
      1 underanvändande
      1 underårig
      3 underarm
      1 underarmarna
      2 underarmen
      1 underarmens
     12 underart
      9 underarten
     13 underarter
      1 underarterna
      1 underater
      1 underavdelning
      1 underavdelningar
      3 underbarn
      3 underben
      4 underbenen
      4 underbenens
      8 underbenet
      1 underbett
      1 underbinda
      1 underblåst
      2 underbyggda
      1 underbyggt
      1 underdelen
      1 underdiagnos
      1 underdiagnosiserat
      1 underdiagnostik
      3 underdiagnostiserat
      1 underdiscipliner
      5 underfamiljen
      1 underfamiljer
      1 underfamiljparvovirinae
      1 underfeminisation
      1 underförstådda
      2 underförstått
      2 underfunktion
      1 underfunktionell
      2 undergå
      1 undergång
      4 undergår
      1 undergick
      1 undergivna
      1 undergörande
      1 undergräva
      9 undergrupp
      7 undergrupper
      1 undergrupperas
      1 undergrupperingar
      1 undergrupperna
      1 underhåll
      1 underhållande
      1 underhållaren
      1 underhållas
      1 underhåller
      1 underhållet
      1 underhållit
      2 underhållning
      1 underhållningssyfte
      2 underhålls
      1 underhållsbehandla
      2 underhållsbehandling
      1 underhållsbehandlingen
      1 underhållsdagar
      1 underhållsdos
      1 underhållsfas
      2 underhållsfasen
      1 underhållsfri
      1 underhållsfunktioner
      1 underhållsmässighet
      1 underhållsmedlen
      1 underhållssäkerhet
      1 underhud
      2 underhuden
      6 underhudsfett
      4 underhudsfettet
      2 underifrån
      1 underjord
      2 underjordiska
      1 underjordsanläggningar
      1 underkäke
      6 underkäken
      2 underkäkens
      1 underkänner
      3 underkant
      1 underkanten
      1 underkastade
      1 underkastar
      1 underkastas
      1 underkastat
      1 underkastelse
      1 underkategoriseras
      1 underkjolar
      4 underkläder
      1 underkläderna
      1 underklädesplagg
      1 underklänning
      2 underklassen
      1 underklasser
      1 underklassificeringar
      4 underklorsyrlighet
      1 underklorsyrlighets
      1 underkonsumtion
      1 underlack
     21 underlag
      8 underlaget
      1 underlägsenhet
      1 underlagskräm
      2 underläkare
      1 underlandet
      4 underläppen
      1 underlåtit
     38 underlätta
      2 underlättade
      1 underlättande
     28 underlättar
     10 underlättas
      1 underlättning
     45 underliggande
      1 underligheter
      2 underligt
      1 underliv
     11 underlivet
      2 underlivets
      1 undermålig
      1 undermaskulinisation
      1 undermedvetna
      7 undernärda
     30 undernäring
      2 undernäringen
      1 undernät
      1 underordnad
      1 underordnade
      1 underordnat
      2 underordning
      3 underordningar
      1 underordningarna
      3 underordningen
      1 underplagg
      4 underproduktion
      1 underpronation
      1 underrapportering
      1 underrätta
      1 underrättad
      1 underrättelseservice
      1 underrättelsetjänster
      1 undersida
     14 undersidan
      1 underskatta
      1 underskattar
      1 underskattats
      1 underskikt
      1 underskötare
      5 undersköterska
      1 undersköterskeprogram
      1 undersköterskeutbildning
      7 undersköterskor
      3 underskott
     69 undersöka
      2 undersökande
      2 undersökandes
      4 undersökaren
      1 undersökarna
     23 undersökas
     17 undersöker
    134 undersökning
     81 undersökningar
      5 undersökningarna
     59 undersökningen
      1 undersökningens
      1 undersöknings
      1 undersökningsgrupp
      1 undersökningsinsatser
      1 undersökningsledare
      3 undersökningsmetod
      1 undersökningsmetoden
      3 undersökningsmetoder
      1 undersökningsmuskeln
      1 undersökningsresultatet
      1 undersökningsteknik
      1 undersökningstid
      1 undersökningstillfälle
      1 undersökningstillfället
     21 undersöks
     11 undersökt
      4 undersökta
      8 undersökte
      3 undersöktes
      6 undersökts
      2 underspecialister
      1 underspecialitet
      2 underspecialiteter
      1 underst
      1 understå
      3 underställd
      1 underställt
      1 understammen
      8 understiger
      1 understimulans
      1 understimulering
      1 understöd
      1 understödd
      1 understöddes
      2 understödjande
      1 understödjas
      1 understryka
      1 understrykas
      1 understryker
      1 understryks
      1 undertill
     10 undertryck
      2 undertrycka
      1 undertryckande
      5 undertrycket
      1 undertrycks
      1 undertrycktes
      1 undertyp
      1 undertyper
      1 underutveckingen
      1 underutvecklad
      1 underutveckling
      1 undervärderar
     11 undervikt
      1 underviktig
      3 undervisa
      3 undervisade
      1 undervisades
      1 undervisar
     13 undervisning
      1 undervisningen
      1 undervisningsämnet
      1 undervisningsinnehåll
      1 underwirebra
      1 undfallenhet
      1 undfly
      2 undgå
      2 undkomma
      1 undkommer
      1 undrar
      1 undrat
      9 undre
      1 undrer
      1 undsätta
      1 undslippa
      1 undulatus
      1 undvara
      2 undvek
      4 undvik
    151 undvika
     13 undvikande
      3 undvikandebeteenden
      2 undvikandet
     18 undvikas
     28 undviker
      1 undvikits
      5 undviks
      1 unesco
     29 ung
     87 unga
      8 ungar
      3 ungarna
      6 ungdom
     57 ungdomar
      4 ungdomarna
      1 ungdomars
      3 ungdomen
      1 ungdomens
      1 ungdomlig
      2 ungdoms
      3 ungdomsåren
      2 ungdomsdiabetes
      1 ungdomsdiabetesinsulinberoende
      1 ungdomsgäng
      3 ungdomsmottagning
      1 ungdomsmottagningar
      1 ungdomsmottagningarna
      1 ungdomspsykiater
      3 ungdomspsykiatrin
      1 ungdomssjukhus
      1 ungdomstid
      8 unge
    287 ungefär
      1 ungefärlig
      3 ungefärliga
      2 ungefärligen
      1 ungeför
      5 ungern
      1 ungerns
      2 ungerska
      1 ungerske
      1 unghundar
      1 ungkarlsliv
      1 ungödlor
      1 ungomen
      2 ungraren
      2 ungt
      1 ungträd
      1 unicef
      1 unicystisk
      2 unie
      1 uniform
      1 uniformer
      1 uniformitet
      7 unik
     10 unika
      2 unikt
     38 unilever
      1 unileverföretagen
      9 unilevers
      2 unilvers
      1 uniokulära
      2 union
      8 unionen
      2 unionens
      4 unipolära
      1 unisonic
      3 unit
      7 united
      1 unity
      1 univ
      1 universalgeniet
      3 universalmedel
      3 universella
      1 universellt
      1 universidad
     74 universitet
      1 universitetcollege
      3 universiteten
      6 universitetet
      1 universitetets
      1 universitets
      1 universitetshögskoleutbildning
      1 universitetsområden
     13 universitetssjukhus
      2 universitetssjukhusen
     18 universitetssjukhuset
      1 universitetssjukhusets
      3 universitetsutbildning
     25 university
     10 universum
      1 unodc
      3 uns
      2 unverdorben
      3 up
      1 upanishaderna
      1 upanishadtraditionerna
      2 upb
      1 upon
    858 upp
     37 uppåt
      1 uppåtbakåtrörelser
      1 uppåtriktad
      1 uppåtstigande
      1 uppåtutåt
      1 uppbåd
      1 uppbär
      1 uppbenbart
      2 uppblandad
      1 uppblandade
      1 uppblåsbar
      1 uppblåsbart
      1 uppblött
      1 uppbromsning
      1 uppbrott
      1 uppbyggande
      1 uppbyggandet
      9 uppbyggd
     16 uppbyggda
     16 uppbyggnad
      5 uppbyggnaden
      5 uppbyggt
      2 uppdagades
      1 uppdagas
      1 uppdagats
      1 uppdal
      1 uppdaterad
      1 uppdaterade
      1 uppdaterades
      1 uppdaterar
      2 uppdateras
      1 uppdaterat
      1 uppdaterats
      1 uppdatering
      3 uppdelad
      1 uppdelade
      6 uppdelas
      2 uppdelat
     13 uppdelning
      1 uppdelningar
      2 uppdelningen
     23 uppdrag
      5 uppdraget
      1 uppdragna
      1 uppdragning
      1 uppdragningskanyl
      1 uppdragningskanylen
      1 uppdragningsskanyl
      1 uppdragsgivare
      2 uppdragsgivaren
      2 uppdragsgivarna
      1 uppdrogs
      1 uppdykande
     19 uppe
      8 uppehåll
      1 uppehälle
      1 uppehåller
      1 uppehållet
      1 uppehållsplatser
      1 uppehållstid
      1 uppehållstidformula
      1 uppehöll
     10 uppemot
      5 uppenbar
      8 uppenbara
      1 uppenbarelse
      5 uppenbarligen
      9 uppenbart
      1 uppfällbar
      1 uppfälld
      1 uppfångade
      5 uppfann
     30 uppfanns
     28 uppfatta
      1 uppfattad
      1 uppfattade
      8 uppfattades
     23 uppfattar
     50 uppfattas
      4 uppfattat
      3 uppfattats
      1 uppfattbarhet
     41 uppfattning
     16 uppfattningar
      3 uppfattningarna
     23 uppfattningen
      2 uppfattningsförmågan
      1 uppfinna
      1 uppfinnandet
      5 uppfinnare
      2 uppfinnaren
      5 uppfinning
      1 uppfinningar
      1 uppfinningen
      1 uppfinningsrikedom
      1 uppflammande
      1 uppfödd
      1 uppfödda
      1 uppfödning
      1 uppfödningen
      1 uppfödningssvårigheter
      3 uppföljande
      1 uppföljd
     20 uppföljning
      3 uppföljningar
      2 uppföljningen
      1 uppföljningsmätningar
      1 uppföljningsstudierna
      3 uppför
      2 uppföranden
     10 uppförandestörning
      1 uppförandestörningar
      2 uppförandet
      1 uppförde
      3 uppfördes
      2 uppförsbacke
      2 uppfostran
      1 uppfräschning
      1 uppfriskande
      2 uppfunnit
      1 uppfunnits
      8 uppfylla
      8 uppfyllas
     11 uppfyllda
      4 uppfyllde
      1 uppfyllelse
     16 uppfyller
      2 uppfylls
      5 uppfyllt
     10 uppgå
      1 uppgående
      9 uppgår
      6 uppgav
      1 uppgavs
      3 uppge
     17 uppger
      3 uppges
      2 uppgett
      5 uppgick
     49 uppgift
      2 uppgiften
     38 uppgifter
      8 uppgifterna
      1 uppgiven
      1 uppgraderades
      1 upphakningar
      1 upphandlades
      1 upphandlingar
      1 upphängda
      1 upphängning
      1 upphängningsanordning
      1 upphävande
      1 upphävandet
      1 upphävda
      1 upphävdes
      1 upphäver
      2 upphävt
      4 upphetsad
      1 upphetsade
      1 upphetsande
     10 upphetsning
      3 upphetsningen
      2 upphetta
      1 upphettad
      2 upphettade
      1 upphettades
      1 upphettar
      5 upphettas
      2 upphettat
      1 upphettats
     15 upphettning
      6 upphöjd
      3 upphöjda
      2 upphöjning
      1 upphöjt
     29 upphör
     13 upphöra
     13 upphörde
     14 upphört
      1 upphostat
      3 upphostning
      2 upphostningar
      1 upphostningarna
    175 upphov
      2 upphovet
      1 upphovsmakare
      2 upphovsman
      1 upphovsmän
      2 uppifrån
      5 uppiggande
      8 uppkallad
      2 uppkallade
      2 uppkallades
      5 uppkallat
      1 uppkallats
      1 uppkastning
      1 uppkastningar
      1 uppklarad
      1 uppklarning
      1 uppknäppta
     17 uppkom
    116 uppkomma
      4 uppkommen
    160 uppkommer
      1 uppkommet
     23 uppkommit
      3 uppkomna
     30 uppkomst
     31 uppkomsten
      1 uppkomstmekanism
      3 uppkomstmekanismer
      1 uppkomstplats
      1 uppköpt
      3 uppl
      1 uppladdningen
      1 uppladdningsbar
      1 uppladdningsbara
      1 upplag
      6 upplaga
      8 upplagan
      2 upplägg
      1 upplägget
      1 uppläggning
      1 upplagor
      1 upplagrade
      1 upplagras
      1 upplagring
      2 uppland
      1 upplandslagen
      2 uppläsningen
     55 uppleva
      1 upplevande
     18 upplevas
      4 upplevd
     14 upplevda
     12 upplevde
      2 upplevdes
     24 upplevelse
      1 upplevelsebaserad
      1 upplevelseliv
     19 upplevelsen
     27 upplevelser
      3 upplevelserna
     98 upplever
     37 upplevs
      8 upplevt
     10 upplösning
      1 upplösningen
      1 upplösningsbara
      1 upplösningsförmåga
      5 upplöst
      2 upplösta
      2 upplöstes
      1 uppluckrad
      1 upplyft
      1 upplyfta
      2 upplyftande
      1 upplyning
      1 upplysas
      1 upplysning
      2 upplysningar
      1 upplysningen
      2 upplysningsmärke
      1 upplysningstiden
      1 upplyst
      4 upplysta
      1 uppmana
      3 uppmanade
      2 uppmanades
      6 uppmanar
      5 uppmanas
      2 uppmanat
      1 uppmanats
      4 uppmaning
      3 uppmaningar
      2 uppmaningen
      6 uppmärksam
     44 uppmärksamhet
      9 uppmärksamheten
      1 uppmärksamhets
      1 uppmärksamhetsalexi
      1 uppmärksamhetsfokus
      1 uppmärksamhetskomponent
      2 uppmärksamhetsstörning
      1 uppmärksamhetsstörningar
      1 uppmärksamhetsstörninghyperaktivitet
     10 uppmärksamma
      3 uppmärksammad
      7 uppmärksammade
      9 uppmärksammades
      1 uppmärksammanden
      2 uppmärksammar
     11 uppmärksammas
      5 uppmärksammat
     11 uppmärksammats
      1 uppmärksamt
      1 uppmärkssamhetssystemet
      2 uppmäta
      1 uppmätande
      1 uppmätbara
      2 uppmätning
      1 uppmäts
      8 uppmätt
      6 uppmätta
      1 uppmättes
      2 uppmätts
      1 uppmjukande
      1 uppmjukas
      1 uppmjukningen
     11 uppmuntra
      1 uppmuntrade
      1 uppmuntrades
      1 uppmuntran
      1 uppmuntrande
      4 uppmuntrar
      2 uppmuntras
     56 uppnå
      3 uppnådd
      4 uppnådda
      2 uppnådde
      1 uppnåddes
      1 uppnåeliga
      1 uppnåeligt
     12 uppnår
     20 uppnås
     11 uppnått
      8 uppnåtts
      1 uppochnedvänt
      1 uppräkning
      1 uppräkningen
      6 upprätt
     11 upprätta
      1 upprättade
      2 upprättades
      3 upprättandet
      1 upprättas
     22 upprätthålla
      2 upprätthållandet
      2 upprätthållas
      1 upprätthåller
      1 upprätthålles
      7 upprätthålls
      1 upprätthölls
      1 upprättstående
      1 uppreglerad
      1 uppreglerade
      2 uppreglerar
      1 uppregleras
      1 uppreglerat
      8 upprepa
      5 upprepad
     44 upprepade
      3 upprepande
      2 upprepar
     13 upprepas
      5 upprepat
      1 upprepats
      4 upprepning
      5 upprepningar
      1 upprepningsbeteende
      1 uppresningslyftar
      1 upprest
      1 uppringarnas
      1 uppritade
      2 uppritningen
      1 upprivna
      1 uppror
      1 upprörd
      3 upprörda
      1 upproret
      1 upprört
      1 upprullningen
     32 uppsala
      1 uppsamla
      1 uppsamlade
      2 uppsamling
      1 uppsamlnigsrör
      2 uppsåt
      1 uppsats
      1 uppsatser
      3 uppsatt
      1 uppsatta
      8 uppsättning
      1 uppsättningar
      3 uppsättningen
      1 uppseende
      3 uppsikt
     15 uppskatta
      5 uppskattad
      5 uppskattade
     10 uppskattar
     24 uppskattas
      6 uppskattat
      2 uppskattats
      4 uppskattning
      7 uppskattningar
      1 uppskattningarna
      2 uppskattningen
     15 uppskattningsvis
      1 uppskjutarbeteende
      1 uppskruvat
      1 uppskurna
      2 uppslagsbok
      2 uppslagsboken
      1 uppslagsord
      1 uppslagsverk
      1 uppslagsverket
      1 uppslukas
     10 uppsöka
      1 uppsökande
      2 uppsökas
      1 uppsöker
      2 uppsöks
      1 uppspänt
      1 uppspelningsmetod
      1 uppsplittrad
    158 uppstå
      1 uppställa
      2 uppställda
      1 uppställde
      3 uppståndelse
    284 uppstår
     38 uppstått
     11 uppstigning
      2 uppstigningar
     29 uppstod
      1 uppstoppad
      1 uppstoppade
      6 uppstötningar
      1 uppsugande
      1 uppsuges
      3 uppsugningsförmåga
      1 uppsugs
      3 uppsvälld
      1 uppsvällda
      2 uppsving
      2 uppsvullnad
      2 uppta
     45 upptäcka
      4 upptäckare
      2 upptäckarna
     14 upptäckas
      8 upptäcker
      1 upptäckresande
     45 upptäcks
     62 upptäckt
      6 upptäckta
     32 upptäckte
     28 upptäckten
     10 upptäckter
      2 upptäckterna
     72 upptäcktes
     11 upptäckts
      1 upptäcktsresor
      1 upptäcktvirussom
     21 upptag
      1 upptaga
      1 upptagande
      8 upptagen
      2 upptagenhet
      9 upptaget
      2 upptagit
      3 upptagna
      4 upptagning
      1 upptagningen
      1 upptagningsmekanism
      1 upptagningsmekanismer
      1 upptagningsvägen
      1 upptänkliga
      6 upptar
     10 upptas
      1 upptecknade
      6 upptill
      1 upptinats
      1 upptining
      1 upptiningsprocessen
      1 upptogs
     48 uppträda
      4 uppträdande
      1 uppträdanden
      1 uppträdandeproblem
      1 uppträdandet
      3 uppträdde
    120 uppträder
      1 upptrappningen
      2 uppträtt
      1 uppväcka
      1 uppväcks
      1 uppväger
      1 uppvaket
      6 uppvaknande
      2 uppvaknanden
      5 uppvaknandet
      4 uppvärmd
      2 uppvärmda
     21 uppvärmning
      1 uppvärmningen
      1 uppvärmningssätt
      3 uppvärmt
      2 uppvätskad
      4 uppväxt
      1 uppväxtår
      2 uppväxtåren
      7 uppväxten
      1 uppväxtförhållanden
      1 uppväxtmiljö
      1 uppväxtvillkor
      1 uppvindar
     15 uppvisa
      1 uppvisade
     59 uppvisar
      3 uppvisas
      5 uppvisat
      1 uppvisningar
      1 uprima
      1 upspel
    265 ur
      1 urakut
      2 uralbergen
      1 urålders
      1 uråldrig
      1 uråldriga
      2 uralit
     32 uran
      1 uranbaserade
      1 uranbrytning
      1 urandioxid
      1 urangult
      1 uranhalter
      1 uranisotoper
      1 uranium
      1 uranockra
      1 uranreserver
      1 uranserien
      1 urantillgångar
      2 urat
      1 uratsten
      2 uratstenar
      2 urban
      1 urbana
      1 urbanae
      1 urbani
      1 urbanisationen
      1 urbaniserade
      1 urbaniseringen
      1 urbefolkningen
      4 urdjur
      6 urea
      1 ureacykeln
      1 ureas
      3 uremi
      1 uretär
      1 uretären
     11 uretrit
      1 urfolksstammar
      2 urgamla
      1 urgammal
      1 urglasförband
      1 urgonaden
      1 urgröpt
      1 uri
      2 uridom
     56 urin
      1 urinanalys
      1 urinavgång
      1 urinbåsan
      2 urinbaserade
      9 urinblåsa
     28 urinblåsan
      1 urinblåsans
      1 urinblåseväggen
      7 urindrivande
      1 urindroppsamlaren
      1 urindroppsamlareuridom
     51 urinen
     15 urinera
      2 urinerade
      2 urinerande
      1 urinerandet
      2 urinerar
     24 urinering
      1 urineringen
      1 urineringens
      4 urinflaska
      3 urinflödet
      1 urinförgiftning
      1 urinfunktioner
      1 uringångarna
      8 urininkontinens
      1 urininkontinenta
      1 urinkateterisering
      2 urinkatetrar
      1 urinkatetrars
      4 urinläckage
      1 urinledande
      1 urinledare
      3 urinledaren
      4 urinledarna
      6 urinmängd
      3 urinmängden
      1 urinmängder
      1 urinmängderna
      1 urinmikroskopi
      1 urinmynning
      1 urinnitriter
      1 urinoarer
      3 urinodling
      1 urinodlingar
      1 urinöret
      1 urinorgan
      1 urinpåsar
      1 urinpåse
      4 urinproduktion
      4 urinproduktionen
      9 urinprov
      3 urinprover
      2 urinretention
      8 urinrör
     33 urinröret
      2 urinrörets
      1 urinrörskatarr
      2 urinrörsmynningen
      1 urinrörsutsöndring
      1 urinsticka
      1 urinsvårigheter
     14 urinsyra
      1 urinsyran
      2 urinträngning
      1 urinuppsamlngspåse
      1 urinutdrivning
      1 urinutsöndring
      1 urinutsöndringen
      5 urinvägar
     18 urinvägarna
      1 urinvägarnas
      1 urinvägen
      3 urinvägs
      1 urinvägsbakterier
      4 urinvägscancer
      1 urinvägshindret
     26 urinvägsinfektion
     26 urinvägsinfektioner
      1 urinvägsinfektionerna
      1 urinvägsorganism
      1 urinvägsproblem
      1 urinvägssjukdom
      1 urinvägssystemet
      1 urinvolymer
      1 urkalkning
      1 urladdas
      1 urladdning
      3 urladdningar
      1 urladdningen
      1 urlaka
      1 urlakade
      1 urlakas
      3 urlakning
      6 urminnes
      1 urnor
      2 urnupna
      7 urografi
      1 urokinas
      3 urolog
      2 urologer
      3 urologi
      1 urologin
      1 urologiska
      1 uroporfyrinogen
      1 urostomi
      1 urringade
      2 urringning
      1 urrivna
      9 ursäkt
     14 urskilja
      2 urskiljas
      1 urskiljde
      1 urskiljer
      1 urskiljs
      1 urskiljtas
      2 urskiljts
      1 urskillning
     80 ursprung
      1 ursprungen
      9 ursprunget
      7 ursprunglig
     40 ursprungliga
      1 ursprungligaste
      1 ursprunglige
     50 ursprungligen
      1 ursprungsbefolkning
      1 ursprungsbetydelse
      2 ursprungscell
      1 ursprungsfärg
      1 ursprungsland
      2 ursprungslandet
      1 ursprungsspänningen
      1 ursprungssubstans
      1 ursprungstumören
      1 ursprungsvävnaden
      1 urt
      1 urta
      1 urtagbar
      2 urtagbara
      2 urti
      1 urtica
      1 urticarial
      3 urtikaria
      1 urtikariatillstånd
      1 urtinktur
      1 uruguay
      2 urushiol
      1 urushioldermatit
     13 urval
      2 urvalet
      1 urvalsgrupp
      1 urvalsgruppen
      1 urvriden
      8 us
    245 usa
      1 usabaserade
      1 usainspirerade
      1 usamriid
     12 usas
      1 usasponsrad
      1 usbanslutning
      1 usc
      3 usd
      2 use
      1 usel
      1 ushers
      1 usk
      2 usp
      1 uspstf
      1 uss
      1 ustilaginomycotina
      1 ustulina
    903 ut
      1 uta
      4 utagerande
      2 utah
    859 utan
      2 utandad
     12 utandning
      8 utandningen
      1 utandningsflöde
      2 utandningsluft
      5 utandningsluften
      1 utandningsprover
      1 utandningsvolym
    103 utanför
      1 utanförroslagstullistockholm
      1 utanförskap
      9 utanpå
      3 utanpåliggande
      2 utarbeta
      1 utarbetad
      5 utarbetade
      2 utarbetades
      1 utarbetande
      1 utarbetar
      1 utarbetas
      3 utarbetat
      6 utarbetats
      1 utarmas
      3 utarmat
      1 utarmats
      9 utåt
      1 utåtgående
      1 utåtledande
      3 utåtriktade
      1 utåtriktat
      6 utbilda
     11 utbildad
     15 utbildade
      1 utbildandet
      4 utbildar
      4 utbildare
      1 utbildaren
      5 utbildas
      4 utbildats
     82 utbildning
      6 utbildningar
      9 utbildningarna
     48 utbildningen
      2 utbildningens
      1 utbildningsform
      2 utbildningskrav
      1 utbildningsnivå
      1 utbildningsnivåer
      1 utbildningsorterna
      1 utbildningsplaner
      1 utbildningsprogrammet
      1 utbildningssyfte
      1 utbildningsträffarna
      1 utblandat
      1 utblåsning
      1 utbölingar
      1 utborrning
      6 utbrändhet
      1 utbreda
     26 utbredd
     15 utbredda
     62 utbredning
      6 utbredningen
     10 utbredningsområde
      1 utbredningsområden
      3 utbredningsområdet
     19 utbrett
      3 utbröt
     64 utbrott
      7 utbrotten
     18 utbrottet
      1 utbrottsfrekvensen
      1 utbrutit
      4 utbudet
      5 utbuktning
      1 utbuktningar
      1 utbyggd
      5 utbyggnad
      1 utbyta
      1 utbytbara
     13 utbyte
      1 utbyter
      2 utbytet
      2 utbytt
      4 utbytta
      1 utc
      1 utdela
      1 utdelades
      5 utdelas
      2 utdelning
      1 utdikning
      1 utdöda
      1 utdömande
      1 utdömas
      3 utdömdes
      1 utdömts
      7 utdragen
      4 utdraget
      4 utdragna
      2 utdragning
      1 utdragningsinstrument
      1 utdrivande
      1 utdrivningsreflex
      1 utdrivningsreflexen
      1 utdrivningsskedet
      1 utdrygning
     18 ute
      2 utebli
     10 uteblir
      7 utebliven
      2 uteblivet
      1 uteblivna
      5 utefter
      1 utelämnade
      1 utelämnades
      1 utepromenader
      1 uterin
      1 uterina
      1 uterintdå
      1 utero
      3 uterus
      1 uteservering
      1 uteserveringar
      1 uteslöt
     26 utesluta
     33 uteslutande
      6 uteslutas
     11 utesluter
      1 uteslutet
      2 uteslutits
      3 utestänga
      2 utestängda
      1 utevistelse
      1 utexaminerade
      1 utexaminerades
      8 utfall
      2 utfaller
      3 utfallet
      5 utfällning
      2 utfällningar
      1 utfälls
      1 utfallsmåtten
      3 utfärda
      1 utfärdad
      5 utfärdade
      2 utfärdades
      5 utfärdar
      3 utfärdas
      5 utfärdat
      1 utfärdats
      1 utfart
      2 utfasning
      3 utflöde
      1 utflödet
      1 utflykter
      1 utflytt
      1 utfodringsförsök
      1 utfodringsstudier
     33 utför
     86 utföra
     12 utförande
      3 utförandeanalys
     12 utföranden
      9 utförandet
      2 utförare
      1 utföraren
      2 utförarna
     58 utföras
     14 utförd
      5 utförda
     11 utförde
     37 utfördes
      1 utföres
      1 utförlig
      1 utförligare
      1 utförligt
      4 utforma
      7 utformad
     12 utformade
      6 utformas
      1 utformat
      6 utformats
     14 utformning
      8 utformningen
    123 utförs
      1 utförsel
      2 utförsgång
      1 utforska
      1 utforskade
      2 utforskande
      1 utforskaren
      1 utforskat
      3 utforskats
      2 utforskning
     10 utfört
      8 utförts
      1 utfrysta
      6 utgå
      5 utgående
     21 utgång
      2 utgången
      1 utgångna
      1 utgångshastighet
      1 utgångsläge
      4 utgångsmaterial
      1 utgångsmaterialet
     11 utgångspunkt
      3 utgångspunkten
      2 utgångspunkter
      1 utgångssättet
     76 utgår
      2 utgått
      2 utgav
      3 utgåva
      5 utgåvan
      2 utgåvor
      5 utgavs
      3 utger
      1 utges
      1 utgett
      4 utgick
      1 utgift
      1 utgifterna
      2 utgivare
      1 utgivaren
      3 utgivna
      1 utgivning
     12 utgjorde
      8 utgjordes
      4 utgjort
      1 utgjorts
      3 utgjutning
    131 utgör
     19 utgöra
      1 utgörande
      5 utgöras
     51 utgörs
      1 utgrävda
      2 utgrävningar
      1 utgrävningarna
      5 uthållighet
      2 uthålligheten
      1 uthållighetsidrott
      2 uthållighetsidrottare
      3 uthållighetsträning
      1 uthärdas
      1 uthyrning
      6 uti
     85 utifrån
      1 utilitaristiskt
      1 utjämna
      1 utjämning
      1 utkämpade
      1 utkanten
      1 utkastform
      1 utkastning
     11 utkom
      2 utkommande
      4 utkommen
      1 utkommit
      1 utkristalliseras
      1 utlakning
      1 utläkningsprocessen
      1 utläkta
      1 utlämnad
      1 utlämning
      1 utländsk
      9 utländska
      1 utlandsresa
      2 utlandsresor
      2 utlåning
      2 utlänningar
      5 utläsa
      1 utlåtande
      1 utlåtanden
      1 utlevelsen
      4 utlöpare
      2 utlopp
      1 utloppet
     23 utlösa
     35 utlösande
      2 utlösare
      1 utlösaren
     18 utlösas
     24 utlöser
     15 utlöses
     10 utlösning
      1 utlösningar
      3 utlösningen
      9 utlöst
      4 utlösta
      1 utlöste
      1 utlösts
      1 utlovade
      1 utlovar
      1 utlyste
      1 utmanade
      3 utmanar
      1 utmanas
      2 utmaning
      6 utmaningar
      1 utmaningarna
      1 utmaningen
      9 utmärkande
      2 utmärkelse
      3 utmärker
      1 utmarkerade
      8 utmärks
      9 utmärkt
      3 utmärkta
      1 utmärkte
      3 utmattad
      8 utmattning
      1 utmattnings
      4 utmattningsbrott
      1 utmattningsdepression
      1 utmattningsfraktur
      1 utmattningssyndrom
      1 utmattningstillstånd
      9 utmed
      1 utmognaden
      1 utmognandet
      3 utmynna
      1 utmynnat
      1 utnämndes
      1 utnämnt
      1 utnämnts
      7 utnyttja
      1 utnyttjad
      1 utnyttjade
      2 utnyttjades
      2 utnyttjande
      1 utnyttjandet
     14 utnyttjar
     19 utnyttjas
      1 utnyttjats
      7 utöka
      3 utökade
      1 utökades
      2 utökas
      2 utökat
     30 utom
      2 utomäktenskapliga
      1 utomäktenskapligt
      1 utomeuropeiska
      8 utomhus
      1 utomhusaktiviteter
      1 utomhusbadande
      2 utomhusvistelse
      2 utomjordingar
      1 utomjordisk
      6 utomkvedshavandeskap
     13 utomlands
      8 utomstående
      1 utöndrar
      1 utopi
      1 utopisk
      1 utopiska
     13 utöva
      3 utövad
      2 utövade
      3 utövades
      5 utövande
      3 utövandet
     23 utövar
      4 utövare
      8 utövaren
      5 utövarna
     12 utövas
      4 utövat
      2 utövats
     64 utöver
      1 utövning
      2 utpekade
      1 utpekar
      1 utpekas
      1 utpetade
      2 utplåna
      1 utplånades
      1 utpmolekyl
      2 utpräglad
      1 utpräglagt
      5 utpräglat
      1 utprovad
      1 utprovade
      1 utprovas
      1 utpumpandet
      1 utpumpning
      1 uträknas
      1 uträkningar
      1 uträkningen
      1 uträtade
      1 uträtat
     17 utreda
      1 utredande
      1 utredare
      2 utredaren
      4 utredarna
      6 utredas
      1 utredd
      4 utredda
      2 utreddes
      3 utreder
     51 utredning
      8 utredningar
      9 utredningen
      1 utredningsmässigt
      1 utredningsmetoder
      1 utredningsresultatet
      2 utreds
      2 utrett
      1 utrikes
      1 utrikespolitik
      8 utröna
      1 utropade
      1 utropat
      1 utropstecken
     16 utrota
      4 utrotad
      4 utrotade
      3 utrotades
      5 utrotas
      2 utrotat
      1 utrötat
      2 utrotats
      4 utrotning
      1 utrotningen
      1 utrotningsförsök
      1 utrotningshotad
      1 utrotningshotade
      1 utrotningskampanj
      1 utrotningsprojekt
      3 utrustad
      8 utrustade
      1 utrustades
      1 utrustat
     34 utrustning
      1 utrustningar
      5 utrustningen
      1 utryckningar
     18 utrymme
      5 utrymmen
      1 utrymmena
      1 utrymmesbesparingar
      1 utrymmesbrist
      1 utrymmeskrävande
      4 utrymmet
      2 utsäde
      1 utsädet
      1 utsågad
      1 utsågades
      1 utsågning
      1 utsago
      1 utsagor
      2 utsägs
      1 utsaltning
      2 utsända
      3 utsänder
      1 utsänt
     11 utsatt
     33 utsatta
      8 utsätta
     14 utsättas
      1 utsatte
     10 utsätter
      7 utsattes
      1 utsatthet
      1 utsattheten
      4 utsättning
      2 utsättningen
     22 utsatts
     57 utsätts
      1 utse
     66 utseende
      1 utseendedefekter
      1 utseendefixering
      1 utseendeförändring
      1 utseendeförändringar
      1 utseendemässiga
      3 utseendemässigt
     22 utseendet
      1 utser
      2 utses
      1 utsetts
      8 utsida
     19 utsidan
      1 utsignalen
      1 utsikten
      1 utsikter
      3 utsikterna
      1 utsirning
      1 utskaffas
      1 utskällde
      1 utskärande
      3 utskärning
      1 utskiljs
      4 utskjutande
     18 utskott
      1 utskrift
      1 utskrivning
      1 utskrivningsprövning
      1 utskuren
      1 utskurna
      1 utsläckta
     49 utslag
     14 utslagen
      4 utslaget
      1 utslagets
      6 utslagna
      1 utslagningsmekanismer
      6 utsläpp
      5 utsläppen
      1 utsläppet
      1 utsläppta
      1 utslätad
      1 utslätning
      1 utslitna
      1 utslocknade
      1 utslungas
      3 utsmyckade
      2 utsmyckning
      1 utsmyckningar
     17 utsöndra
      1 utsöndrad
      3 utsöndrade
      1 utsöndrades
      2 utsöndrande
     42 utsöndrar
     70 utsöndras
      2 utsöndrat
      2 utsöndrats
      1 utsöndrig
     29 utsöndring
      4 utsöndringar
     24 utsöndringen
      1 utsöndringens
      1 utsot
      1 utsövd
      7 utspädd
      4 utspädda
      3 utspädning
      1 utspädningar
      3 utspädningen
      1 utspädningsfaktorn
      1 utspärrade
      2 utspätt
      2 utspelar
      2 utspridda
      1 utsprutas
      4 utstå
      3 utstående
      1 utställd
      3 utställning
      2 utställningen
      1 utställningskuvöserna
      1 utstjälpningar
      1 utstötas
      1 utstötningsprocesser
      2 utstötta
      1 utsträcker
     79 utsträckning
      1 utsträckningar
      1 utsträckt
      1 utsträckte
      1 utstrålad
      1 utströmmar
      1 utströmning
      1 utströmningen
      1 utsvettning
      1 uttag
      1 uttaga
      1 uttaget
      1 uttagna
      1 uttagning
      1 uttagningshjälp
     10 uttal
      2 uttala
     12 uttalad
     15 uttalade
      3 uttalande
      2 uttalanden
      2 uttalandet
      3 uttalar
     13 uttalas
      8 uttalat
      1 uttalats
      9 uttalet
      1 uttalsavvikelser
      1 uttalsförändring
      1 uttalsförändringar
      1 uttalsträning
      1 uttalsutvecklingen
      2 uttänjda
      1 uttänjning
      1 uttolkningen
      1 uttömda
      1 uttömmande
      4 uttömning
      3 uttömningar
      2 uttömningen
      2 uttorkad
      2 uttorkade
      3 uttorkande
     30 uttorkning
      1 uttorkningstillstånd
      2 utträde
      2 uttråkad
      1 uttröttade
      1 uttröttande
     83 uttryck
     10 uttrycka
      5 uttryckas
     10 uttrycken
     14 uttrycker
     32 uttrycket
      3 uttryckligen
      1 uttryckligt
      9 uttrycks
      1 uttrycksförmågan
      3 uttrycksformer
      1 uttrycksfullt
      1 uttryckslöst
      9 uttryckt
      5 uttryckte
      1 uttryckts
      1 uttsatts
      1 uttycket
      1 uttyckt
      2 uturkroppenupplevelse
      1 utvädring
      3 utväg
      2 utvägen
      3 utvald
      4 utvalda
      1 utvalt
      1 utvanns
      4 utvärdera
      1 utvärderad
      2 utvärderade
      3 utvärderades
      6 utvärderar
      3 utvärderas
      3 utvärderat
      3 utvärderats
     36 utvärdering
      6 utvärderingar
      1 utvärderingen
      1 utvärderings
      1 utvärderingsbart
      7 utvärtes
      1 utvärtesparasit
      1 utväxling
      2 utväxt
      1 utväxta
      1 utväxter
    104 utveckla
     20 utvecklad
     69 utvecklade
     75 utvecklades
      1 utvecklande
      9 utvecklandet
     87 utvecklar
      1 utvecklaren
      1 utvecklarna
    188 utvecklas
     43 utvecklat
     69 utvecklats
    148 utveckling
      1 utvecklingan
      2 utvecklingar
    101 utvecklingen
      3 utvecklingens
      1 utvecklingrubbningar
      1 utvecklingsbana
      1 utvecklingsbar
      1 utvecklingsbetingad
      1 utvecklingsbetingade
      1 utvecklingscentret
      1 utvecklingsdefekt
      1 utvecklingsdyslexi
      2 utvecklingsfasen
      1 utvecklingsfaser
      1 utvecklingsgången
      1 utvecklingshistoria
      1 utvecklingskedjan
      1 utvecklingskedjor
     20 utvecklingsländer
      9 utvecklingsländerna
      1 utvecklingsländernade
      1 utvecklingslära
      1 utvecklingslinje
      1 utvecklingsmässiga
      3 utvecklingsnivå
      1 utvecklingsnivåer
      1 utvecklingsperioden
      1 utvecklingsprocessen
      2 utvecklingsprojekt
      1 utvecklingspsykiatri
      3 utvecklingspsykologi
      1 utvecklingspsykologiskt
      4 utvecklingsrubbning
      1 utvecklingssamarbete
      1 utvecklingssjukdomarna
      1 utvecklingsstadier
      1 utvecklingsstadium
      3 utvecklingsstörda
      1 utvecklingsstördas
     59 utvecklingsstörning
      4 utvecklingsstörningar
      1 utvecklingsteam
      1 utvecklingsteorierna
      1 utvecklingstillstånd
      3 utvidga
      2 utvidgad
      6 utvidgade
      5 utvidgar
      7 utvidgas
      2 utvidgat
      1 utvidgats
     10 utvidgning
      1 utvidgningen
      1 utvilad
      6 utvinna
      6 utvinnas
      5 utvinner
      3 utvinning
     13 utvinns
      2 utvisa
      1 utvunnen
      1 utvunnet
      2 utvunnit
      3 utvunnits
      1 uuh
      5 uv
      6 uva
      1 uvabehandling
      1 uvabsorberare
      1 uvacrispa
      2 uvåg
      1 uvbestrålning
      1 uvea
      1 uveit
      1 uvfilter
      9 uvi
      2 uvier
      2 uvisymptom
      1 uvlampor
      7 uvljus
      1 uvs
      3 uvskydd
      1 uvskyddet
      1 uvstrålar
      3 uvstrålning
      1 uvulopalatopharyngoplastik
      1 uysal
      1 u�z
      1 uzbekistan
     19 v
      1 vaayu
      1 väbel
      1 väblar
      2 vacca
    107 vaccin
     45 vaccination
      7 vaccinationen
      5 vaccinationer
      2 vaccinationerna
      2 vaccinationsgrad
      1 vaccinationsgraden
      1 vaccinationskampanjer
      1 vaccinationsmetoden
      7 vaccinationsprogram
      3 vaccinationsprogrammet
      1 vaccinationsprogrammets
      1 vaccinationstillfället
      1 vaccine
     13 vacciner
     11 vaccinera
      4 vaccinerad
     18 vaccinerade
      1 vaccinerande
      1 vaccinerar
     13 vaccineras
      3 vaccinerats
     11 vaccinering
      1 vaccineringsgrad
      2 vaccinerna
     37 vaccinet
      1 vaccinforskning
      1 vaccinforskningen
      1 vacciniavirus
      1 vaccinimmunitet
      1 vaccinrelaterad
      1 vaccinsäkerhet
      1 vaccinutveckling
     11 väcka
      1 väckande
      2 väckarklocka
      1 väckas
      4 vacker
      9 väcker
      4 vackert
      1 väckningshjälpmedel
      9 vackra
      1 vackrare
      1 vackraste
      7 väcks
      1 väckt
      6 väckte
      2 väcktes
      1 väckts
      1 vacuum
    327 vad
      5 vådabekämpning
      1 vådabeskjutning
      1 vadderad
      1 vadderade
      1 vadderat
      4 vaddering
     18 väder
      4 väderförhållanden
      2 väderkartor
      2 väderlek
      1 väderleken
      3 vaderna
      1 väderspänningar
      1 väderstreck
      2 vädjan
      1 vädjar
      1 vädjat
      1 vadlånga
      1 vadmuskeln
      1 vadmuskelpumpen
      1 vadmuskulaturen
      1 vadomfång
      2 vädra
      3 vädras
      3 vädret
      2 vadstena
      3 vag
      7 våg
     53 väg
      8 vaga
      1 våga
      7 väga
      2 vagabond
      1 vågade
      2 vägande
      1 vågar
     27 vägar
      1 vägarbetare
      1 vägarbetaren
      3 vägarbete
      2 vägarbeten
      2 vagare
      3 vägarna
      1 vägbanor
      1 vägbara
      2 vägbeläggning
      1 vägbeläggningen
      1 vagbhata
      1 vagbhatas
      1 vägbulan
      1 vägbulor
      1 vägbulors
      3 vägde
      1 vågdeformationens
      1 vågen
     41 vägen
     23 väger
      1 vägförhållanden
      1 vågformen
      5 vågformer
      9 vägg
      1 vagga
      2 vaggar
     18 väggar
      5 väggarna
      1 väggbeklädnad
      7 väggen
     27 vägglöss
     10 vägglössen
      6 vägglus
      1 vägglusarter
      1 vägglusavföring
      1 vägglusbekämpning
      1 vägglusdrabbad
      1 vägglusdrabbat
     35 vägglusen
      7 vägglusens
      2 vägglusfälla
      1 vägglushona
      1 vägglushonan
      1 väggluspopulationen
      1 vägglusproblemet
      1 vägglussanering
      1 vägglussaneringar
      1 vägglussläktet
      1 vägglusspår
      1 vaggningen
      1 väggplattor
      1 väggrepp
      2 vägguttaget
      1 väghållaren
      1 vågig
      2 vågiga
     20 vagina
      1 vaginae
     12 vaginal
     10 vaginala
      1 vaginalinlägg
     14 vaginalis
      1 vaginalpessar
      1 vaginalring
      2 vaginalringar
      1 vaginalringen
      1 vaginalsex
     10 vaginalt
     10 vaginan
      1 vaginans
      1 vaginata
      8 vaginism
      2 vägkant
      1 vägkanten
      2 vägkanter
      5 vägkorsning
      2 vägkorsningen
      2 väglag
      5 våglängd
      1 väglängd
      1 våglängden
      4 våglängder
      1 våglängderna
      1 våglängdsområden
      1 våglängdsområdet
      4 vägleda
      2 vägledande
      1 vägledd
      1 vägledda
      1 vägleder
      6 vägledning
      2 vägledningen
      5 vägmärken
      1 vägmärkena
      1 vägmärket
      1 vågmönster
      1 vagnar
      1 vagnberga
      1 vagnhärad
      3 vägningsfilter
      1 vägojämnheter
      1 vägområden
     12 vågor
      2 vågorna
      6 vägrade
      8 vägrar
      3 vägrat
      2 vågrätt
      3 vägrenar
      2 vågrörelse
      1 vågrörelseperiod
      3 vägs
      1 vägsalt
      1 vägskatetrar
      2 vägt
      1 vägtrafikdefinitioner
      2 vagus
      1 vagusnerven
      1 vägverkets
      1 väja
      3 väjningsplikt
      1 väjningspliktsmärken
      9 vaken
     14 vakenhet
      2 vakenheten
      1 vakenhetgrad
      1 vakenhets
      4 vakenhetsgrad
      1 vakenhetsgraden
      1 vakenhetshöjande
      1 vakenhetssänkt
      1 vakenhetsstörningar
      4 vakenhetsterapi
      3 vakenhetsterapin
      1 vakenhetsterapins
      7 vaket
     17 vakna
     14 vaknar
      1 vaknat
      2 vaksam
      1 vaksamhet
      1 vaksamheten
      1 vaksamma
      1 vakt
      3 väktare
      1 väktarutbildade
      1 vaktas
      1 vaktbolag
      1 vaktel
      1 vaktkapten
      1 vaktkår
      2 vakuol
      5 vakuum
      1 vakuumaspirering
      1 vakuumextirpation
      1 vakuumförpackningar
      1 vakuumpannor
      1 vakuumpump
      2 vakuumrör
      2 vakuumsalt
      2 vakuumsystem
     29 val
     99 väl
      1 valaciclovir
      1 valaciklovir
      2 välanpassade
      1 valar
      2 välavgränsade
      1 välbärgade
     21 välbefinnande
      6 välbefinnandet
      1 välbegåvade
      1 välbehag
      1 välbehagskänsla
      4 valben
      1 valbens
      1 välbeprovad
      1 valbo
      1 vald
     37 våld
      3 valda
      9 valde
      1 väldefinierat
      1 valdes
      1 väldet
    112 väldigt
      4 väldoftande
      1 väldokumenterad
      1 väldokumenterade
      2 väldokumenterat
      1 väldokumunterat
      1 väldränerad
      1 väldränerade
      1 vålds
      1 våldsam
      1 våldsamhetsrisk
      9 våldsamma
      1 våldsammare
      4 våldsamt
      1 våldsanvändning
      1 våldsbenägna
      8 våldsbrott
      1 våldsbrotten
      1 våldsbrottslingar
      1 våldshämmande
      2 våldsmonopol
      1 våldsmonopolet
      1 våldsutbrott
      1 våldsutövare
      1 våldsutövning
     10 våldtäkt
      1 våldtäkter
      1 våldtäktsman
      1 våldtäktsmannen
      1 valegnani
      2 valen
      2 valens
      1 valensbindningsteori
      1 valenseffekten
      1 valenselektroner
      1 valenselektronerna
      1 valensen
      2 valent
      1 valentindagsmassakern
      9 valet
      1 väletablerad
      2 väletablerade
      3 välfärd
      1 välfärden
      1 välfärdsproblem
      1 välfärdsstaten
      1 välfärdsstatens
      2 valfiskben
      1 välförgrenad
      1 välformad
      1 valfri
      2 valfrihet
      1 valfriheten
      6 valfritt
      1 valfunktionärer
      1 valfusk
      1 välgång
      1 valgiserande
      3 välgjorda
      1 välgjort
      1 välgörande
      1 välgöraren
      1 valgum
      1 validera
      1 validitet
      1 valin
      1 välinformerad
     42 välja
      5 väljas
     30 väljer
      8 väljs
      4 välkänd
     15 välkända
      1 välkändhet
      6 välkänt
      2 valkar
      2 valkas
      2 valkning
      4 välkomna
      1 valla
      1 vålla
      1 vållade
      2 vållande
      1 vallar
      3 vållar
      1 vållat
      1 vallatae
      1 vållats
      1 vallebona
      3 vallentin
      1 valleskog
      1 vällevnadssjukdomarna
      1 vallfärdade
      1 vallfärden
      1 vallfärder
      1 vallhundar
      1 välling
      1 vällingen
      1 vallmosaft
      1 vallmotorp
      3 vallmoväxter
      1 vallo
      1 vällovliga
      1 vällukt
      9 välmående
      1 välmåga
      1 välnärda
      1 valnöt
      1 valnötslik
      2 valnötter
      1 valobservatörer
      2 valpar
      1 valpat
      1 välplanerad
      1 valproat
      1 valproater
      1 valproatsyndrom
      5 valproinsyra
      4 valpsjuka
      2 valpsjukevirus
      1 välrenommerad
      1 välrenommerade
      1 valresultat
      2 valresultatet
      1 valrossben
      1 valsar
      1 välsigna
      1 välsignelse
      1 välsmakande
      1 valspråk
      1 välstånd
      1 välstuderade
      1 valsverket
      6 valt
      1 valtaktik
      1 vältränad
      4 vältränade
      1 valtrex
      1 valts
      1 välts
      1 valujev
      4 valuta
      1 valutaförordningen
      1 valutakod
      1 valutalagen
      1 valutan
      3 valutareserv
      2 valutavärde
      1 välutförda
      2 välutvecklad
      1 välutvecklade
      3 välutvecklat
      1 valvbåge
      1 välvd
      1 välvda
      1 valvet
      1 valvsena
      2 våmmen
      1 vampyrattribut
      1 vampyrism
      1 vampyrsjukan
     17 van
      4 vän
     10 vana
      4 vanan
      1 vanartig
      2 vancomycin
      2 vancomycinresistenta
      2 vänd
      6 vända
      1 vandalism
      2 vändas
      6 vände
     10 vänder
      1 vändning
     11 vandra
      3 vandrande
     17 vandrar
      4 vandrat
      1 vandring
      1 vandringssägen
      1 vandringsspindel
      2 vänds
      1 vanebildande
      1 vanemässig
      4 vanemässiga
      1 vanemässigt
      1 vanemönster
      1 vänersborg
      1 vanessa
      2 vanestörningar
      1 vanför
      9 vanföreställning
     73 vanföreställningar
     15 vanföreställningarna
      3 vanföreställningen
      1 vanföreställningsdiagnos
      1 vanföreställningsstörningar
     24 vanföreställningssyndrom
      1 vanföreställningssyndromen
      1 vanföreställningssynrom
      1 vanföreställningsyndrom
      1 vanförställningen
      1 vanhedra
      1 vaniljkräm
      1 vaniljsås
      1 vaniottii
      3 vänja
      3 vänjer
      5 vankomycin
    256 vanlig
      2 vänlig
    291 vanliga
      2 vänliga
    151 vanligare
    125 vanligast
    364 vanligaste
      1 vanlige
    425 vanligen
    443 vanligt
      1 vänligt
    290 vanligtvis
      8 vann
     21 vänner
      2 vänners
      8 vanor
      1 vanorna
      1 vanprydande
      1 vanquin
      1 väns
      5 vansinne
      1 vansinnesköra
      2 vänskap
      1 vänskapen
      1 vänskapliga
      1 vänskapsrelationer
      1 vansköta
      2 vanställande
      2 vanställda
      2 vanställningar
     75 vänster
      1 vänsterform
      1 vänsterförmaksförstoring
      1 vänsterhandtaget
      1 vänsterhänt
      2 vänsterhänta
      2 vänsterkammare
      1 vänsterkammaren
      1 vänsterradikala
      1 vänsterradikaler
      1 vänstersidig
      2 vänstersidiga
      1 vänstersidigt
      8 vänstertrafik
      1 vänstertrafiken
      1 vänstervarianterna
      1 vänstervridna
     35 vänstra
      2 vant
      1 vänt
     12 vänta
      3 väntade
      3 väntan
      1 väntande
      1 vantar
      8 väntar
      2 väntas
      1 väntat
      1 vänterhjärtat
      2 väntetid
      1 väntetiden
      1 vantolkas
      1 vantolkningar
      1 vantro
      1 väntrum
      4 vanvård
     48 vapen
      1 vapenbärare
      1 vapendragare
      1 vapenindustrin
      1 vapenlås
      1 vapenlicens
      1 vapenlicenser
      2 vapenplutonium
      2 vapenskåp
      1 vapenskölden
      1 vapenställ
      3 vapensystem
      1 vapentekniska
      1 vapentyper
      2 väpnade
      1 väpnat
      3 vapnen
      7 vapnet
      3 vapnets
      3 vaporizer
      1 vaporizern
   1501 var
     52 vår
   1793 vara
     27 våra
      7 varade
      1 varadenguefebern
      1 varaivärldenvaro
      6 varaktig
      6 varaktiga
     19 varaktighet
      2 varaktigheten
      8 varaktigt
      3 varan
      1 varanarter
      2 varande
    137 varandra
      6 varandras
      8 varanen
      5 varanens
      7 varaner
      3 varanerna
     11 varannan
      1 varannat
      1 varanödlans
      1 varansamlingar
      8 varanus
     35 varar
      1 vårarna
      1 vårärt
      5 varat
      1 varatt
     71 varav
      1 varbakterier
      1 varberg
      3 varbildning
      1 vårblomma
      2 varböld
      1 vårby
      1 vårbyfittjatrakten
    129 vård
     16 värd
      3 vårda
      3 värda
      3 vårdades
      7 vardag
     12 vardagen
      4 vardaglig
     21 vardagliga
      4 vardagligare
     16 vardagligt
      2 vardags
      1 vardagsaktiviteter
      1 vardagsanvändning
      1 vardagsliv
      1 vardagslivet
      1 vardagsnära
      1 vardagsplagg
      1 vardagspsykopat
      2 vardagspsykopaten
      1 vardagssammanhang
      1 vardagssjukvården
      2 vardagsspråk
      3 vardagsspråket
      1 vardagstal
      1 vårdalternativ
      3 vårdande
      1 vårdanstalterna
      2 vårdar
      1 värdar
      1 vårdaren
      1 vårdarens
      1 värdarter
     10 vårdas
      2 vårdat
      3 vårdats
      1 vårdavdelning
      3 vårdavdelningar
      1 vårdavtal
      1 vårdbehovet
      1 vårdberoende
      2 vårdbiträden
      1 vårdbundet
      3 värdcell
      7 värdcellen
      2 värdcellens
      9 vårdcentral
      4 vårdcentralen
      7 vårdcentraler
      5 vårdcentralerna
      1 vårdcentralernas
      9 värddjur
      2 värddjuren
      4 värddjurens
      4 värddjuret
      2 värddjurets
     42 värde
      7 värdefull
      3 värdefulla
      1 värdefullare
      3 värdefullt
      1 värdeladdade
      1 värdeladdning
      1 värdelös
      3 värdelösa
      1 värdelöst
     50 vården
     96 värden
      6 värdena
      3 vårdens
      6 värdens
      1 värdepappersform
     15 vardera
      5 värdera
      1 värderad
      1 värderade
      1 värderades
      1 värderar
      2 värderas
      5 värdering
      7 värderingar
      1 värderingen
      1 värderingsförändringar
      2 värderingstabell
      4 värdesätta
      2 värdesätter
     24 värdet
      1 värdeteoretiska
      1 värdeteori
      1 vårdformen
      1 vårdformer
      1 vårdfrågor
      6 vårdgivare
      1 vårdgivaren
      1 vårdgivarna
      1 vårdguiden
      1 vardguidense
      4 vårdhem
      6 vårdhund
      2 vårdhundar
      3 vårdhunden
      1 vårdhundens
      1 vårdhundshundsföraren
      1 vårdhundsprojekt
      1 vårdhygien
      1 vårdhygieniska
      1 vårdidealen
      4 värdighet
      2 värdigt
      3 vårdinrättningar
      2 vårdinsatser
      1 vårdinstitutioner
      1 vårdkontakten
      1 vårdkvalitet
      1 vårdlinjen
      1 vårdmiljö
      3 värdmödraskap
      1 vårdnadsfrågor
      2 vårdnivå
      2 vårdområdet
      3 värdorganism
      3 värdorganismen
      4 värdorganismens
      1 vårdpedagogik
     14 vårdpersonal
      4 vårdpersonalen
      1 vårdpersonals
      2 vårdplatser
      1 vårdprofessionell
      1 vårdrelaterad
      3 vårdrelaterade
      1 värdskap
      1 vårdslöshet
      1 värdspecificitet
      1 värdspecifika
      1 vårdsystemen
      1 vårdsystemets
      2 vårdtagare
      3 vårdtid
      1 vårdtider
      1 vårdtillfällen
      1 vårdutbildning
      2 värdväxt
      2 värdväxten
      3 värdväxtens
      4 vårdvetenskap
      1 vårdyrken
     64 vare
     24 varefter
     10 varelse
     11 varelsen
      1 varelsens
     12 varelser
      4 varelses
     30 våren
      1 varenda
      1 vareniklin
      3 varet
    110 varför
      2 varfyllda
     12 varg
      1 vargangrepp
      9 vargar
      7 vargen
      1 varghund
      1 vargjägare
      1 varglever
      3 vargliknande
      1 vargref
      1 vargsopp
      1 vargspindlar
      1 vargunge
      2 varhärd
      1 varhärden
      3 vari
      7 variabel
      2 variabelt
      1 variabilis
      2 variability
      3 variabla
      3 variabler
      2 varians
     69 variant
     22 varianten
     90 varianter
      8 varianterna
     21 variation
      4 variationen
     17 variationer
      5 variationerna
      1 varibeln
      7 varicella
      2 varicer
     63 variera
      1 varierad
     10 varierade
     47 varierande
    156 varierar
      3 varieras
      7 varierat
      1 varietéer
      3 varieteter
     13 varifrån
      2 varig
      3 variga
     12 varigenom
      2 varigt
     45 varilux
      1 variluxglaset
      1 varinnehållet
      4 variola
      1 variolavirus
     12 variolisation
      1 variolisera
      2 variolisering
    254 varit
      2 varius
      2 varixblödning
      2 värja
    254 varje
     35 värk
      1 värka
      2 värkande
      1 värkarbete
      1 värkarbetet
     37 varken
      7 värken
      3 värktabletter
      1 värktabletterna
      1 vårlandskapet
      5 värld
      6 världar
      1 världarna
    247 världen
      1 världenden
     71 världens
      1 världensamhällena
      2 världs
      2 världsaidsdagen
      1 världsaidskampanjen
      1 världsallergiorganisationen
      3 världsalltet
      1 världsandens
      1 världsbefolkningen
      2 världsbild
      1 världscancerdag
      1 världscancerdeklaration
      1 världscancerkongresser
      4 världsdelar
      1 världsdelarna
      1 världsfrälsare
      1 världsgrunden
      2 världshälsodagen
     39 världshälsoorganisationen
      8 världshälsoorganisationens
      1 världshälsoorganistionen
      1 världshälsorapporten
      1 världshärskare
      2 världshaven
      1 världshistorien
      1 världshistoriens
      1 världsjälen
      1 världskongress
     46 världskriget
      4 världskrigets
      1 världsledande
      1 världslepradagen
      1 världsliga
      1 världslivsmedelsprogrammet
      1 världsmusik
      1 världsomfattande
      1 världsorganisation
      1 världspremiären
      1 världsprincip
      1 världsproblem
      1 världsproduktionen
      1 världspsykiatriförbundet
      1 världsserien
      3 världssjälen
      1 världssvälten
      1 världsträd
      1 världsträdet
      1 världsutsällningen
      2 världsvida
      1 världsvitt
      1 varligt
      1 vårlökssläktet
     14 varm
     23 varma
      7 värma
      1 värmanordning
      6 varmare
      2 värmas
      2 varmaste
      1 varmblodig
      6 varmblodiga
      2 värmdes
     38 värme
      1 värmebehandla
      1 värmebehandlad
      1 värmebehandlade
      1 värmebehandlas
      3 värmebehandling
      1 värmebölja
      1 värmeböljor
     11 varmed
      2 värmedesinfektion
      2 värmedyna
      3 värmedynor
      1 värmeelement
      1 värmefiltar
      1 värmeförluster
      1 värmegrad
      2 värmeisolerande
      1 värmeisolering
      3 värmekällan
      3 värmekänsliga
      1 värmekänsligt
      2 värmekollaps
      1 värmekramper
      1 värmekuddar
      2 värmekudde
      1 värmelampa
      1 värmeledningen
     11 värmen
      2 värmeödem
      4 värmeökning
      1 värmepanna
      1 värmepannor
      1 värmeplåster
      1 värmeproducerande
      1 värmepumpar
      1 värmer
      3 värmerelaterade
      1 värmesäng
     14 värmeslag
      1 värmeslaget
      1 värmetåligt
      1 värmetorkskåp
      1 värmeutslag
      1 värmeutstrålning
      1 värmeuttag
      1 värmeuttagen
      1 värmeutvecklingen
      2 värmevallning
      1 värmevallningar
      5 värmland
      1 värmlands
      2 varmluft
      1 varmmangel
      1 varmpressning
      1 varmrökt
      1 varmrökta
     12 värms
      1 värmslag
     29 varmt
      1 varmtkallt
      1 vårmusseron
      1 vårmusseronen
      3 varmvatten
      1 varmvattenanslutna
      1 varmvattenbassäng
      1 varmvattenrör
      1 varmvattenrören
      1 varmvattensystemet
      5 varna
      2 varnade
     39 varnar
      2 varnas
      6 varning
      6 varningar
      1 varningsfilm
      1 varningslista
      2 varningsmärke
      9 varningsmärken
      1 varningsmärket
      5 varningssignal
      1 varningssignaler
      1 varningsskylt
      1 varningsskyltar
      1 varningsskylten
      4 varningstecken
      1 varningstecknen
      3 varningstext
      4 varningstexter
      1 värnplikt
      2 värnplikten
      2 värnpliktiga
     11 varor
      2 varorna
      1 varorsakat
     13 varpå
      1 värphöns
     17 värre
    104 vars
      1 varsam
      1 varsamhet
      2 varsamt
      1 vårsäsongen
      1 varse
      1 varsebli
      6 varseblivning
      1 varseblivningarna
      1 varseblivningen
      3 varseblivningshjälpmedel
      1 varsin
      1 vårskotten
      8 värst
     36 värsta
      2 vårstädning
     19 vart
     18 vårt
      9 värt
      2 vårta
      1 vårtan
      4 vartannat
      1 vartdera
      2 vårtecken
      3 vartefter
      5 vårtgård
      4 vårtgårdar
      1 vårtgårdarna
      6 vårtgården
      1 vårtig
      1 vårtiga
      1 vårtlika
      9 vårtor
      5 vårtorna
      1 vårtsvin
      4 varulexikon
      2 varulv
      1 varum
      5 varumärke
      7 varumärken
      1 varumärkena
      1 varumärkeslöftet
      9 varumärket
      7 varunamn
      5 varunamnet
      1 varunder
      1 varunummer
      7 varv
      1 varva
      1 varvar
      3 varvas
      1 varvätska
      1 varvet
     57 varvid
      1 varvsarbetare
      1 varvsindustrin
      2 vas
      1 vasa
      1 väsa
      5 väsande
      1 vasco
      1 vascular
      1 vasculosa
      1 vasektomi
      1 vasektomier
      4 vaselin
      1 vaseline
      1 vasen
     11 väsen
      1 väsenet
      1 väsenskilda
      1 väsensskild
      4 väsentlig
      2 väsentliga
      1 väsentligaste
      4 väsentligen
      1 väsentlighet
     15 väsentligt
      2 vaser
      1 vask
      4 väska
      1 väskan
      6 vaskulär
      5 vaskulära
      1 vaskulärdemens
      6 vaskulit
      1 vaskuliter
      1 vaskulitsjukdomar
      3 väsningar
      2 vasoaktiva
      3 vasodilatation
      1 vasogent
      1 vasokonstrikterande
      4 vasokonstriktion
      1 vasokonstriktionen
      1 vasokonstriktor
      2 vasomotorcentrum
      9 vasopressin
      1 vasopressinadh
      1 vasopressinbalansen
      1 vasospasm
      1 vasospasmen
      1 vass
      4 vassa
      1 vasslen
      1 vassopresin
      2 vasst
      1 vasstrån
     15 väst
      8 västafrika
      3 västafrikanska
      1 västar
      3 väster
      3 västerås
      3 västerbotten
      2 västerbottens
      2 västergötland
      8 västerlandet
      1 västerlandets
     10 västerländsk
     27 västerländska
      1 västerländskt
      2 västerlänningar
      1 västerneran
      1 västernorrlands
      5 västerut
      4 västeuropa
      1 västeuropeiska
      4 västindien
      1 västjylland
      4 västkust
      2 västkusten
      1 västkustskolan
      3 västländer
      1 västländerna
      1 västlig
      2 västliga
      1 västmanland
      2 västmanlands
     21 västra
      1 västsverige
     47 västvärlden
      1 västvärldens
      1 västvärldspiercing
      1 våt
      1 vata
      3 våta
      1 våtare
      1 våtbastu
      2 våtbastun
      2 våtdräkt
      2 väte
      2 väteatom
      2 väteatomen
      2 väteatomerna
      1 vätebinder
      6 vätebindningar
      1 vätebindningarna
      1 vätebromid
      6 vätecyanid
      1 vätefluorid
      1 vätejon
      6 vätejoner
      1 vätejonkoncentrationen
      1 vätejonkoncentrationerna
      2 vätekarbonat
      1 vätekarbonatjoner
      5 väteklorid
      1 väteorganeller
     34 väteperoxid
      1 väteperoxidens
      1 väteperoxidnedbrytande
      2 väteperoxidsalva
      1 vateri
      2 vätesuperoxid
      6 vätgas
      1 vätgasen
      1 våthet
      1 våtmarker
      1 våtmarksbiotoper
      1 våtmarksmygga
      1 våtplåtar
      1 våtrakning
    153 vätska
     31 vätskan
      1 vätskans
      1 vätskatarmsaft
      2 vätske
      1 vätskeabsorberande
      1 vätskeadministrering
      7 vätskeansamling
      1 vätskeansamlingar
      1 vätskeavstötande
      5 vätskebalans
      4 vätskebalansen
      2 vätskebehandling
      8 vätskebrist
      1 vätskebristen
      5 vätskedrivande
     14 vätskeersättning
      1 vätskeförande
      1 vätskeförlust
      3 vätskeförlusten
      1 vätskeförluster
      1 vätskeförlusterna
      1 vätskeformiga
      4 vätskefylld
      4 vätskefyllda
      1 vätskehalten
      7 vätskeintag
      2 vätskeintaget
      1 vätskekontroll
      1 vätskekromatografi
      2 vätskeläckage
      1 vätskeläckaget
      1 vätskelik
      2 vätskemängden
      1 vätskenivån
      1 vätskeöverbelastning
      1 vätskereabsorption
      1 vätskestygn
      1 vätskesvullen
      5 vätsketillförsel
      1 vätsketrycket
      1 vätskeuppbyggnaden
      3 vätskeutgjutning
      1 vätskeutträde
      1 vätskevandring
     22 vätskor
      6 vätskorna
      3 vått
    360 vatten
      4 vattenånga
      2 vattenansamlingar
      1 vattenanvändning
      1 vattenavstötande
      1 vattenbalansen
      2 vattenbaserade
      3 vattenbaserat
      2 vattenbehållare
      2 vattenbehandlingen
      1 vattenbindande
      1 vattenblandning
      1 vattenborttagande
      1 vattenbråck
      1 vattenbrist
      1 vattenbufflar
      2 vattenburen
      1 vattenbyten
      1 vattendensiteten
      1 vattendirektivet
     10 vattendrag
      1 vattendragen
      1 vattenekvivalenta
      1 vattenfärger
      1 vattenfast
     14 vattenförgiftning
      1 vattenförgiftningen
      1 vattenföroreningar
      1 vattenförvaltning
      3 vattenfri
      1 vattenfria
      1 vattenfylld
      1 vattenfyllda
      1 vattenfylls
      1 vattenfyllt
      1 vattengående
      1 vattenglas
      1 vattengränser
      2 vattenhål
      1 vattenhalten
      1 vattenhaltig
      1 vattenhastighet
      1 vattenhastigheter
      1 vattenhjulet
      1 vatteninhållande
      1 vatteninnehållet
      1 vattenintag
      1 vattenkar
      3 vattenkastning
      1 vattenklar
      1 vattenklosetter
      1 vattenklosetternas
      1 vattenkoncentrationen
      1 vattenkoppor
      1 vattenkranarna
      1 vattenkvalitet
      1 vattenlandning
      1 vattenlås
      3 vattenledningar
      1 vattenledningsnätet
      2 vattenledningssystem
      7 vattenlevande
      1 vattenlinjen
      1 vattenliv
      1 vattenlöpning
      4 vattenlösliga
      1 vattenlöslighet
      9 vattenlösligt
      9 vattenlösning
      2 vattenlösningar
      1 vattenlösningen
      1 vattenmängden
      1 vattenmetabolism
      1 vattenmiljö
      1 vattenmiljöer
      1 vattenmiljön
      4 vattenmolekyler
      1 vattenmyndigheten
      1 vattennät
      1 vattennäten
      1 vattennivån
      1 vattenorganismer
      2 vattenpipan
      5 vattenpipor
      1 vattenpolitiska
      1 vattenpump
      1 vattenpumpen
      1 vattenrelaterat
      4 vattenrening
      2 vattenreningsverk
      2 vattenrör
      1 vattensamling
      3 vattensamlingar
      1 vattensilver
      7 vattenskalle
      1 vattenskräck
      1 vattensnäcka
      1 vattensystem
      1 vattentankar
      2 vattentemperatur
      1 vattentemperaturer
      1 vattenterapins
      1 vattentryck
      2 vattentunn
      1 vattenutsöndring
      1 vattenväxter
      1 vattenväxters
      8 vattenytan
      1 vattenytans
      2 vattenytor
      1 vättern
      1 vätterns
     20 vattkoppor
      2 vattkoppsinfektion
      2 vattnas
      3 vattnen
     75 vattnet
      2 vattnets
      2 vattnig
      1 vattniga
      1 vattnigare
      2 vattnigt
      2 vattuskräck
      1 vattusot
      1 vaumesle
      1 vauquelin
      1 vävd
      1 vävda
      1 vävde
      1 väven
    100 vävnad
     48 vävnaden
      2 vävnadens
     92 vävnader
     32 vävnaderna
      1 vävnaders
      2 vävnads
      1 vävnadsarkitektur
      1 vävnadsbehov
      2 vävnadsbildning
      1 vävnadsbitar
      1 vävnadsbrist
      2 vävnadsceller
      1 vävnadsdestruktion
      3 vävnadsdöd
      1 vävnadsdonation
      1 vävnadsdoppler
      3 vävnadsfaktor
      1 vävnadsförändring
      2 vävnadsförändringar
      1 vävnadsförändringen
      1 vävnadsformer
      1 vävnadsförstoring
      1 vävnadshypoxi
      2 vävnadslager
      1 vävnadslagren
      1 vävnadslevande
      1 vävnadslim
      1 vävnadslimmet
      1 vävnadsodling
      1 vävnadsökning
     11 vävnadsprov
      7 vävnadsprover
      1 vävnadsprovet
      1 vävnadsprovets
      2 vävnadsreaktion
      1 vävnadsreaktioner
      5 vävnadsskada
      1 vävnadsskadliga
      5 vävnadsskador
      1 vävnadsskikt
      1 vävnadssmärta
      1 vävnadsspecifika
      1 vävnadstillväxt
      1 vävnadstryck
      1 vävnadstyper
      1 vävnadsundergång
      1 vävnadsutrymmet
      1 vävnadsvänliga
      2 vävnadsvätska
      1 vävnadsvätskan
      4 vax
      1 vaxa
     48 växa
      2 vaxad
     12 växande
      1 växandet
      2 vaxartad
      1 vaxas
      1 vaxat
      1 växel
      3 växelspänning
      2 växelström
      1 växelvarma
      6 växelvis
      1 vaxer
    117 växer
      1 vaxet
      5 växla
      3 växlande
      6 växlar
      3 växlat
      1 växlingar
      8 vaxning
      1 vaxningen
      1 vaxprodukter
      1 vaxpropp
      1 vaxproppar
     45 växt
      1 växtämnen
      1 växtantioxidanter
      3 växtart
      3 växtarter
      2 växtätare
      1 växtätares
      1 växtbekämpningsmedel
      1 växtbetingelserna
      3 växtdelar
      1 växtdödande
     13 växte
      1 växtembryot
     81 växten
     11 växtens
     97 växter
     10 växterna
      6 växternas
      4 växters
      1 växtextrakt
      2 växtfamilj
      1 växtfärger
      1 växtfärgning
      1 växtförhållanden
      1 växtförökning
      1 växtgiftintoxikationer
      1 växtgrupper
      1 växthormoner
      1 växthuseffekten
      1 växthusgas
      2 växthusgaser
      1 växthusgaserna
      1 växtinnehållet
      1 växtkemist
      1 växtkropp
      1 växtlighet
      1 växtlokaler
      1 växtmaterial
      1 växtmöjligheter
      1 växtnamn
      1 växtöstrogener
      1 växtplats
      1 växtplatser
      3 växtriket
      1 växtsaft
      4 växtsaften
      1 växtsäsong
      5 växtsätt
      1 växtsättet
      3 växtsjukdom
      1 växtsjukdomar
      2 växtskyddsmedel
     17 växtsläkte
      1 växtsläktet
      1 växtsorter
      1 växtvärk
      1 vbatteri
      1 vc
      1 vcr
      2 vd
      1 vdrl
      8 veck
     71 vecka
      1 veckad
      4 veckade
     33 veckan
      2 veckans
      1 veckar
      4 veckas
      1 vecken
      1 vecklar
      1 veckning
      1 vecko
      1 veckodagarna
    179 veckor
     11 veckorna
     10 veckors
      1 vector
      1 vectorerna
      8 ved
      3 veda
      1 vedaratade
      1 vedartad
      1 vedartade
      3 vedaskrifterna
      1 vedeldad
      1 vedeldade
      3 veden
      1 vedens
      6 vederbörande
      2 vederbörandes
      1 vederbörligt
      6 vedertagen
      4 vedertaget
      8 vedertagna
      4 vediska
      1 vedrester
      1 veer
      8 vegan
     22 veganer
      1 veganföreningen
      4 veganism
      1 veganismen
      1 vegankost
      1 veganrörelsen
      8 vegansk
      2 veganska
      1 vegas
      1 vegasautomaterna
      1 vegetabiler
      1 vegetabilia
      9 vegetabilisk
      4 vegetabiliska
      2 vegetabiliskt
     11 vegetarian
     14 vegetarianer
      1 vegetarianerna
      4 vegetarianism
      3 vegetarianismen
      8 vegetarisk
      3 vegetariska
      1 vegetariskt
      3 vegetation
      1 vegetationen
      1 vegetationsrika
      2 vegetativt
      1 vegf
      1 vehicle
      1 veil
      1 veitsdansen
      1 veitstanz
      2 veka
      1 vekar
      1 vektor
      3 vektorburen
      2 vektorer
      1 vektorn
      1 vektorskop
      4 velat
      1 velofarynx
      1 velokardiofacialt
      1 velum
     19 vem
     11 ven
      9 vena
      1 venae
      2 venedig
      1 venedigs
      5 venen
      1 venens
     38 vener
      1 venereal
      3 venereolog
      1 venereologen
      1 venereologer
      1 venereologmottagningar
      2 veneriska
     18 venerna
      1 venerologimottagningar
      1 venesectio
      1 venet
      1 venetiansk
      1 venetianskorna
      1 venetianskt
      1 venetus
      2 venezuela
      6 venkateter
      1 venkatetern
      2 venkatetrar
      1 venklaffar
      1 venlafaxin
      2 venoler
      2 venolerna
      1 venom
      4 venoocklusiv
     10 venös
      9 venösa
      8 venöst
      1 venosus
      1 vensonografi
      1 vensystem
      1 vensystemet
      4 ventil
     21 ventilation
      4 ventilationen
      2 ventilationsanläggningar
      1 ventilationsförmågan
      1 ventilationshål
      2 ventilationskanaler
      1 ventilator
      1 ventilatorassocierad
      1 ventiler
      1 ventilera
      1 ventilerad
      2 ventileras
      1 ventilering
      1 ventoline
      1 ventrala
      1 ventriculi
      1 ventriculus
      1 ventrikelcancer
      1 ventrikelfladder
      8 ventrikelflimmer
      1 ventrikelinnehåll
      1 ventrikellumen
      2 ventrikeln
      1 ventrikelområdet
      4 ventrikelsköljning
      2 ventrikelsköljningen
      1 ventrikelsond
      1 ventrikelsystem
      3 ventrikelsystemet
      1 ventrikeltakykardi
      2 ventriklar
      3 ventriklarna
      1 ventrikulära
      1 ventrikulografin
     18 ventrombos
      1 ventrombosen
      1 ventromediala
      1 ventryck
      1 ventrycket
      1 venusfigurerna
      1 venusgördel
      1 venuskrona
      1 venväg
      1 vepor
      1 vepser
      2 vera
      1 veran
      2 verapamil
      1 veraphamil
      1 veratrum
      3 verb
     10 verbal
      4 verbala
      1 verbalamnesi
      5 verbalt
      5 verbet
      1 verbform
      1 verbformen
      1 verdurins
      3 verifiera
      2 verifierad
      1 verifierade
      1 verifieras
      2 verifierat
      1 verifierbara
      1 verifiering
      1 verint
      1 verizon
     16 verk
     38 verka
     11 verkade
     72 verkan
      8 verkande
    176 verkar
      2 verken
     20 verket
      3 verkets
      7 verklig
     17 verkliga
     23 verkligen
      5 verklighet
     44 verkligheten
      2 verklighetens
      1 verkligheter
      1 verklighets
      1 verklighetsförädnring
      1 verklighetsfrämmande
      1 verklighetsnivån
      6 verklighetsuppfattning
      3 verklighetsuppfattningen
      6 verkligt
      1 verkning
      7 verkningar
      1 verkningarna
      2 verkningsgrad
      1 verkningsgraden
      2 verkningslös
      3 verkningslösa
      8 verkningsmekanism
      5 verkningsmekanismen
      3 verkningsmekanismer
      1 verkningsmekansim
      1 verkningsprofil
      1 verkningssätt
      1 verkningssättet
      2 verkningstid
     15 verksam
     58 verksamhet
     23 verksamheten
      1 verksamhetens
      9 verksamheter
      1 verksamheterna
      1 verksamhetsbeteckning
      1 verksamhetschef
      3 verksamhetsfält
      2 verksamhetsfälten
      2 verksamhetsområde
      1 verksamhetsområdet
      1 verksamhetstillsyn
     34 verksamma
      1 verksammare
     14 verksamt
      1 verkstad
      1 verkstadsindustrin
      3 verkställa
      6 verkställande
      1 verkställandet
      1 verkställde
      1 verkställdes
      1 verkställigheten
      1 verkställs
      1 verkställts
     28 verktyg
      2 verktygen
      1 verktyget
      1 vermicularis
      4 vermiformis
      3 vermikulit
      1 vermox
      1 verner
      2 vernon
      1 vernus
      1 verrucosa
      1 vers
      5 versa
      2 versailles
      1 versaler
      1 versicolor
      4 version
     15 versionen
      3 versioner
      1 versionerna
      1 versraderna
      2 versus
      1 vertebrae
      1 vertebrater
      1 verticalis
      1 vertigo
      9 vertikal
      6 vertikala
      1 vertikalare
      4 vertikalt
      1 verum
      3 very
      1 vesaas
      2 vesalius
      3 vesica
      1 vesicarius
      1 vesicula
      3 vesikel
      1 vesikelexocytosen
      1 vesikeln
      5 vesiklar
      1 vesiklarna
      1 vesikouretär
      2 vesikulär
      1 vestibularisdelen
      1 vestibularmembranet
      1 vestibuli
     12 vestibulit
      1 vestibulitis
      1 vestibulitsyndrom
      1 vestibulocochlearis
      1 vestibulum
      1 vestitus
     56 vet
     21 veta
      1 vetande
      1 vetandet
      7 vete
      2 veteallergi
      1 vetegroddsolja
      1 vetemjöl
     23 vetenskap
     21 vetenskapen
      2 vetenskapens
      3 vetenskaper
     31 vetenskaplig
    103 vetenskapliga
     54 vetenskapligt
      1 vetenskapsakademien
      1 vetenskapsakademiens
      1 vetenskapsexperter
      2 vetenskapsgren
      4 vetenskapsmän
      3 vetenskapsmannen
      1 vetenskapsmännen
      1 vetenskapsområde
      1 vetenskapspris
      2 vetenskapsrådet
      1 vetenskapsteori
      1 veteproteinet
      1 veteraner
      7 veterinär
      1 veterinära
      1 veterinärassistenter
      3 veterinären
      8 veterinärer
      1 veterinärförbund
      1 veterinärhomeopati
      1 veterinärintyg
     10 veterinärmedicin
      1 veterinärmedicine
      9 veterinärmedicinen
      1 veterinärmedicinsk
      5 veterinärmedicinska
      1 veterinärmottagnningar
      1 veterinärpraktiker
      1 veterinärstudenter
      1 veterinärvård
      1 veterinäryrket
      1 vetskap
      1 vetskapen
      2 vetter
      1 vettigare
      2 vev
      1 vevade
      2 vevar
      1 vf
      1 vformade
      1 vhs
    150 vi
    377 via
      5 viagra
      1 vialarter
      1 vialer
      1 vialsläktet
      1 viau
      8 vibration
     10 vibrationer
      1 vibrationsangioödemet
      1 vibrationsgivare
      1 vibrationsskada
      1 vibrationsskador
      2 vibrator
      1 vibratorer
      1 vibrera
      2 vibrerande
      4 vibrerar
      1 vibrio
      6 vice
      1 vickande
      2 vickrar
      1 vicks
      1 vicryl
      3 victor
      3 victoria
   3372 vid
     22 vida
    219 vidare
      1 vidarebefordrar
      1 vidarebefordras
      1 vidaredistribueras
      1 vidarekopplade
      1 vidareoxidation
      2 vidareutbilda
      1 vidareutbildade
      1 vidareutbildas
      4 vidareutbildning
      1 vidareutbildningar
      1 vidareutveckla
      1 vidareutvecklade
      2 vidareutvecklades
      2 vidareutvecklas
      1 vidareutvecklat
      3 vidareutveckling
      1 vidarkliniken
      1 vidast
      1 vidd
      2 videgård
      1 videgårds
      5 video
      1 videoexempel
      1 videokonferensutrustning
      1 videomaterial
      2 videosignaler
      1 videsläktet
      1 vidfästningsredskap
      3 vidga
      6 vidgade
      1 vidgades
      1 vidgande
      6 vidgar
     10 vidgas
      2 vidgats
      4 vidgning
      1 vidgningens
      1 vidhäftad
      1 vidhålla
      1 vidhåller
      2 vidmakthålla
      1 vidmakthållandet
      5 vidmakthåller
      3 vidmakthålls
      1 vidrigt
      1 vidrör
      2 vidröra
      1 vidrörning
      2 vidrört
      3 vidskepelse
      1 vidskepelsen
      1 vidskepliga
      1 vidsynta
     13 vidta
      1 vidtaga
      1 vidtagits
      1 vidtagna
      2 vidtar
      5 vidtas
      1 vidtillgänglig
      3 vidtog
      1 vidvinkelseendet
      6 vietnam
      1 vietnamkriget
      3 viewpoint
      2 vifta
      1 viftar
      3 vigd
      1 vigeland
      2 vigilans
      1 vigiles
      2 vigneaud
      1 vigselböcker
      1 vihta
      8 vii
      9 viii
      1 viiis
      1 vijar
      8 vika
      2 vikas
      1 viken
      3 viker
      1 viking
      1 vikingarna
      1 vikingatid
      2 vikingatiden
      1 vikitiga
      1 vikningen
      2 viks
     89 vikt
      1 viktad
      1 viktbaserad
     21 vikten
      1 vikter
      1 viktförändring
      1 viktförändringar
      2 viktförlust
      1 vikthållning
    142 viktig
    100 viktiga
     12 viktigare
      3 viktigast
     91 viktigaste
    234 viktigt
      1 viktimologin
      2 viktkontroll
      1 viktminskade
      2 viktminskande
     20 viktminskning
      3 viktminskningen
      1 viktminskningsfas
      1 viktminskningsfasen
      1 viktminskningsmetod
      1 viktminskningsmetoder
     21 viktnedgång
      1 viktningsfaktor
      7 viktökning
      1 viktor
      2 viktoria
      1 viktorianska
      1 viktorias
      1 viktprocent
      2 viktprogram
      1 viktprogrammet
      1 viktunderhållande
      8 viktuppgång
      1 vikunja
      1 vil
     51 vila
      1 vilade
      1 vilan
      9 vilande
     11 vilar
      1 vilat
      2 vilcabamba
      5 vild
     20 vilda
      1 vilden
      2 vildformen
      1 vildkanin
      1 vildmarken
      2 vildpersilja
      5 vildsvin
      1 vildsvinet
      1 vildsvinshår
      3 vildväxande
     33 vilja
     22 viljan
      1 viljande
      1 viljans
      1 viljeansträngning
      1 viljehandlingar
      1 viljeliv
      4 viljelivet
      2 viljelös
     11 viljelöshet
      2 viljelösheten
      2 viljemässiga
      2 viljemässigt
      2 viljestyrd
      6 viljestyrda
      1 viljestyrt
      1 viljor
    336 vilka
     12 vilkas
    255 vilken
   1364 vilket
      1 vilketvilka
    397 vill
      1 villa
      1 villafastighetsförsäkring
      1 village
      1 villahem
      1 villarpaskott
      1 villbär
     18 ville
      1 villebråd
      1 villefranche
      1 villekunde
      1 villfarelse
      1 villfarelser
      6 villi
      3 villiga
      1 villighet
     22 villkor
      1 villkorad
      1 villkoras
      2 villkoren
      1 villus
      2 villusatrofi
      1 viloekg
      2 vilohem
      1 vilohjärtfrekvensen
      2 vilomembranpotential
      1 vilomembranpotentialen
      1 viloperioder
      1 vilopotential
      1 vilopotentialen
      2 vilopuls
      2 vilosmärta
      1 viloställen
      1 vilotiden
      1 vilotillståndet
      3 vilseledande
      1 vilseleder
      1 vilstadium
     17 vilt
      1 viltfaunan
     17 vin
      6 vinäger
      1 vinägeraktig
      1 vinbär
      1 vinbärsblad
      1 vinbärsgelé
      1 vinbergssnäckan
      1 vinbergssnäckor
      1 vince
      2 vincent
      1 vincentius
      1 vincenz
      4 vinci
     11 vind
      3 vindar
      1 vindblommiga
      1 vindblommor
      1 vindburna
      8 vinden
      1 vindförhållanden
      2 vindpollinerade
      1 vindpustar
      1 vindriktningen
      1 vindrutan
      3 vindruvor
      1 vinealis
      5 viner
      1 vinexporten
      9 vingar
      1 vingård
      1 vingarna
      1 vingelsjuka
      1 vingkantade
      1 vinglister
      2 vinglösa
      1 vingpenna
      1 vinka
      8 vinkel
      1 vinkelkoordinater
      1 vinkelmätare
      2 vinkeln
      2 vinkelräta
      1 vinkla
      1 vinklad
      1 vinklade
      6 vinklar
      3 vinklingen
      1 vinkristin
      4 vinna
      1 vinnare
      4 vinner
      2 vinning
      1 vinningen
      1 vinningens
      1 vinruta
      4 vinst
      1 vinsten
      3 vinster
      1 vinsterna
      1 vinstgivande
      1 vinstintressen
      1 vinstpotential
      4 vinter
      1 vinterdäck
      1 vinterdepressioner
      1 vinterdräkt
      1 vinterfjäll
      1 vinterförhållanden
      4 vintergäck
      1 vintergäcken
      1 vintergäckssläktet
      2 vintergrön
      1 vintergröna
      2 vinterhalvåret
      4 vinterkräksjuka
      1 vinterkräksjukan
      1 vinterkriget
      1 vintermånaderna
     20 vintern
      1 vintersötesläktet
      1 vintertid
      1 vintrarna
      1 vintyper
      1 vinyasayoga
      2 vinylklorid
      1 violence
      4 violett
      6 violetta
      1 violfärgad
      1 violletleduc
      2 vioxx
      2 vipeholm
      1 vipeholms
      2 vipeholmsexperimenten
      1 vipeholmstoffee
      1 vipeholmsundersökningarna
      1 viper
      1 vipera
      1 viperida
      1 vippärt
      1 virade
     20 viral
      4 virala
      2 viralt
      1 virar
      3 virchow
      1 virginal
      1 virginala
      5 virginia
      1 virginiana
      1 virginiatobaken
      1 viridansstreptocker
      1 virilisation
      2 viriliserande
      1 virilisering
      1 virion
      6 virke
      2 virket
      1 virologi
      1 virologisk
      2 vironerna
      2 virosa
      2 virtual
      6 virtuell
      4 virtuella
      1 virtuellt
      4 virulens
      1 virulensen
      3 virulent
    190 virus
      1 virusämnet
      1 virusbakterier
     10 virusen
      1 virusens
      1 viruses
    137 viruset
     12 virusets
      2 virusfamilj
      1 virusfamiljen
      1 virusförekomsten
      1 virusgenomet
      1 virushalten
      4 virushepatit
      1 virushepatiter
     10 virusinfektion
      2 virusinfektionen
     11 virusinfektioner
      1 virusisolatet
      1 virusisolation
      1 virusisolering
      1 virusisoleringstesterna
      1 virusmängden
      4 virusnivåer
      1 virusnivåerna
      1 virusorsakad
      2 virusorsakade
      1 viruspartikelns
      5 viruspartiklar
      2 viruspartiklarna
      6 viruspneumoni
      1 viruspneumonier
      1 virusprotein
      1 virusproteinernas
      2 virusproteinet
      1 virusreplikation
      1 virusrna
      9 virussjukdom
      3 virussjukdomar
      1 virussjukdomarna
      1 virussjukdomen
      1 virussorterna
      1 virusspecifik
      1 virusspridning
      1 virusspridningen
      4 virusstammar
      2 virusstammen
      1 virustammar
      1 virustyp
      2 virustyper
      1 virusvektorer
      1 virvel
      1 virvelavlossningar
     47 vis
     85 visa
      3 visad
    114 visade
     12 visades
      1 visan
    251 visar
     23 visas
    215 visat
     20 visats
      1 visavi
      1 visby
      3 visceral
      1 viscerala
      1 visdom
      1 visdomständer
      1 visdomständerna
      3 viset
      1 vishnudevananda
      2 vision
      1 visionärt
      2 visionen
      3 visioner
      1 visitkort
      1 viska
      1 viskade
      1 viskande
      1 viskar
      4 viskeralt
      1 viskningar
      2 viskositet
      1 viskositeten
      2 visköst
      1 vismutgallat
      1 vismutnitrat
      1 visningsenhet
      1 vison
      1 vispgrädde
    249 viss
   1031 vissa
      1 visselpipor
     14 visserligen
      1 vissheten
      1 vissla
      1 vissnade
      1 vissnar
      1 vissnat
     73 visst
      6 visste
      1 vistades
     23 vistas
      1 vistats
      4 vistelse
      1 vistelsen
      1 vistelser
      3 visualisera
      1 visualiserar
      3 visualisering
      7 visuell
     13 visuella
      1 visuellspatial
      1 visumkrav
      1 visuospatiala
      4 visus
     61 vit
    119 vita
      1 vitae
      6 vitaktig
      1 vitaktiga
      3 vital
     12 vitala
      5 vitalism
      2 vitalismen
      1 vitalismens
      1 vitalistisk
      1 vitalistiska
      1 vitalitetshormon
      4 vitalkapacitet
      4 vitalkapaciteten
      1 vitalparametrar
     45 vitamin
      2 vitaminbrist
      1 vitamind
      1 vitaminen
     28 vitaminer
      2 vitaminerna
      1 vitaminet
      1 vitamintillskott
      2 vitare
      1 vitblommande
      1 vite
      1 vitfärgning
      1 vitglödning
      3 vitgörande
      1 vitgröe
      1 vitgröna
      1 vitgula
      2 viti
     16 vitiligo
      1 vitiligoforskning
      1 vitium
      7 vitlök
      1 vitoxel
      1 vitreus
      1 vitrifikation
      1 vitro
      1 vitrofertilisering
      2 vitröta
      1 vitryssland
      1 vitsäpel
      1 vitsäper
      5 vitsippa
      5 vitsippan
      1 vitsippans
      1 vitsipporna
     28 vitt
      1 vittene
      3 vittnar
      5 vittnen
      1 vittnesmål
      1 vittnesmålet
      2 vittnesuppgifter
      1 vittvätt
      2 vitus
      1 vitvara
      1 vitvaruföretaget
      1 vivax
      1 vivekananda
      1 vivian
      1 vivipara
      2 vivisektion
      2 vivotif
      2 vivus
      2 vkorc
      1 vkts
      1 vlaardingen
      4 vlcd
      2 vlciak
      2 vlcsfa
      1 vlsi
      1 vm
      1 vmd
      2 vocalise
      2 vocalismuskeln
      2 vocalisutskotten
      1 voice
      1 voipkommunikation
      1 vokabulär
      1 vokabulären
      1 vokal
      1 vokala
      1 vokalen
      7 vokaler
      3 vokalerna
      2 vokalernas
      2 vokalis
      1 vokalklanger
      1 vokalligamentet
      2 vokalliknande
      1 vokalljud
      3 vol
      1 volantes
      3 volfram
      1 volframjodiden
      1 volframmetall
      1 volgasvamp
      3 volt
      1 voltaire
      1 voltaren
      1 voltdiv
      1 voltmeter
      1 voltmetrar
      1 voltruta
      1 volts
      1 voluma
      1 volume
      1 voluminös
      6 voluntarism
      2 voluntarismen
      1 voluntarismens
      1 voluntas
      4 voluven
      1 volvere
      3 volvulus
     31 volym
      1 volymelement
     18 volymen
      1 volymenhet
      6 volymer
      1 volymförändring
      1 volymkontrollerad
      1 volymprocent
      1 volymreceptorer
      1 volyms
      2 volymstyrd
      1 volymsubstitution
      1 volymtidsenhet
      1 vomeronasala
      1 vomiting
      1 vomitoria
     39 von
      1 voodoo
      1 vördas
      2 vördnadsvärde
     11 vore
      1 voriconazol
      1 voro
      1 vortexflödesmätaren
      1 vot
      2 voxel
      1 voxlarna
      1 voyager
      4 voyeurism
      1 vpt
      1 vrår
      3 vre
      3 vred
      1 vredesutbrott
      1 vredet
      1 vreds
      1 vreinfektion
      1 vretyp
      2 vrickning
     11 vrida
      1 vridas
      2 vridbar
      4 vrider
      1 vridit
      3 vridna
      1 vridningsaxeln
      1 vridningsbenägna
      1 vrids
      5 vridspoleinstrument
      1 vrist
      1 vs
      1 vu
      1 vulgär
      1 vulgära
      2 vulgaris
      1 vulgärnamnet
      1 vulkaner
      1 vulkanisering
      1 vulkaniseringen
      1 vulkaniseringsprocessen
      1 vulkanisk
      1 vulkanutbrott
      1 vulkningstemperatur
      5 vulva
      1 vulvan
      1 vulvapapillomatos
      1 vulvärt
      1 vulvavestibulit
      2 vulvodyni
      1 vulvovestibulit
      6 vunnit
     65 vuxen
      1 vuxenåldern
      1 vuxenåren
      1 vuxenblöjor
      1 vuxendöv
      2 vuxendöva
      1 vuxenhabilitering
      1 vuxenincest
      2 vuxenliv
      3 vuxenlivet
      1 vuxenpsykiater
      2 vuxenpsykiatrin
      1 vuxenrollen
      1 vuxenutbildningen
      1 vuxenvärlden
      8 vuxit
    237 vuxna
      1 vuxnarisken
      1 vuxnas
      2 vuxne
      1 vuxnes
      2 vv
      1 vvs
      1 vvsinstallatörer
      2 vy
      1 vyer
      1 vyplastik
      2 vzv
      1 vzvvaccination
      8 w
      2 waal
      1 waalskrafterna
      1 waardenburgs
      1 wadegiles
      1 wae
      2 waerland
      1 waerlandianer
      1 wägner
      2 wagnerjauregg
      1 wahlbom
      1 wahlöös
      1 wahn
      1 wahwah
      1 wahwaheffekt
      1 wais
      1 waistestet
      1 waisthipratio
      1 wakame
      2 wake
      5 wakefield
      5 waksman
      1 waldenström
      1 waldenströms
      1 waldorfpedagogiken
      1 waldorfpedagogikens
      1 waldorfskolorna
      2 wales
      1 walker
      1 wallmark
      2 wälöfwande
      9 walter
      1 wang
      1 waorani
      2 waran
      8 warfarin
      1 warfarinresistens
      1 warming
      1 warner
      1 warrant
      3 warranter
      1 wartec
      1 was
      3 washington
      2 washkansky
      1 wassermannreaktion
      2 water
      1 �watereri
      1 watergate
      1 waterhousefriderichsens
      4 watson
      1 watts
      1 wavefront
      1 waves
      1 wawawa
      2 way
      1 ways
      1 wdr
      1 web
      1 webb
      1 webbbaserat
      1 webben
      7 webbplats
      1 webbplatsen
      4 webbplatser
      1 webmd
      1 websiter
      2 websterstratton
      1 wechsler
      2 wechslers
      1 wechslertest
      1 wechslertesten
      1 wegeners
      1 wehrmacht
      1 weichselbaum
      1 weigelts
      1 weils
      1 weimartiden
      5 weiss
      1 weizmanninstitutet
      1 wellbeing
      7 wells
      1 weltschmerz
      1 wensman
      1 wentin
      1 were
      1 werner
      9 werners
      4 wernickes
      2 werther
      1 werthereffekt
      1 werthers
      6 west
      1 wester
      1 westergren
      1 westermani
      4 western
      1 westling
      1 westlund
      1 westminster
      1 wfot
     19 wfp
      4 wfps
      1 wg
      1 wha
      2 what
      1 when
      3 whiplash
      1 whiplashkommission
      1 whiplashkommissionen
      1 whiplashpatienter
      2 whiplashrelaterade
      1 whiplashskada
      1 whiplashskadade
      2 whiplashskador
      1 whiplashtrauma
      1 whiplashvåld
      1 whipples
      1 whitei
      2 whitening
     72 who
      1 wholaboratorier
      1 whoprojekt
      1 whoregioner
     22 whos
      1 whoskalan
      2 whr
      1 whytt
      1 wichita
      1 wid
      3 wide
      1 widerström
      1 wieloch
      6 wien
      1 wieröe
      1 wiesel
      1 wifalk
      1 wiggers
      1 wiggersdiagrammet
      1 wigmore
      2 wikipedias
      2 wilde
      1 wilder
      2 wilderness
     11 wilhelm
      1 wilkens
      1 wilkins
      1 willans
      1 willebrandfaktorn
      3 willebrands
      2 willem
      1 willemkarel
     27 william
      1 williams
      1 willibald
      1 willis
      1 willumsen
      1 wilms
      1 wilson
      1 wilsonii
      2 wilsons
      1 wimbledonmästerskapen
      1 winchester
      1 winnicott
      1 winter
      1 wirzjustice
      1 wisborg
      1 wisconsin
      1 wisconsinmadison
      9 with
      1 witten
      2 wittenoom
      2 wkromosom
      2 wöhler
      1 wolbachia
      1 wolffchaikoffs
      2 wolffparkinsonwhitesyndromet
      1 wolffska
      2 wolfgang
      1 wolo
      1 wolves
      2 womens
      1 wonderbra
      1 wonderful
      1 woodward
      1 woody
      1 workers
      2 working
      1 works
      1 workshop
     10 world
      1 worlds
      1 woronowii
      1 wortley
      1 wounds
      1 wps
      2 wpwsyndrom
      4 wpwsyndromet
      1 wrestlern
      1 wrestling
      2 wretlind
      1 wrist
      1 writebol
      3 wuchereria
      1 würzburg
      1 wuul
      4 ww
      1 wwwclinicaltrialsgov
      1 wwwinfomedicase
      1 wwwsosse
      1 wwwzumbacom
      1 wyeomyia
      3 wyeth
     26 x
      1 xantenses
      1 xanthoderma
      1 xanti
      1 xantinalkaloid
      1 xantinförgiftning
      1 xantomatos
      1 xaser
      1 xau
      1 xaxeln
      1 xbenthet
      1 xcm
      8 xenobiotika
      5 xenon
      1 xenoöstrogen
      1 xenoöstrogener
      2 xenopsylla
      1 xenos
      2 xenotransplantation
      1 xeomin
      1 xerosis
      1 xerostomi
      1 xhtml
      1 xi
      3 xii
      2 xiii
      1 xiis
      1 ximeng
      1 xiv
      5 xkromosom
      4 xkromosomen
      1 xkromosomer
      1 xml
      1 xochimilco
      1 xolotl
      1 xplattorna
      1 xpotenser
      1 xray
      1 xskalan
      1 xv
      1 xx
      2 xxxviii
      1 xyfoster
      1 xygenotyp
      2 xykromosomer
      1 xylentoluen
      1 xylocaininjektion
      1 xylos
      1 xyoscilloskop
      6 xyy
      5 xyymän
      1 xyypojkar
      1 xyysyndrom
      6 y
      1 yakaspråket
      1 yakuzans
      5 yang
      1 yanomamostammens
      1 yasargilfrån
      1 yasser
      4 yaws
      1 yaxeln
      1 year
      1 yemen
      1 yerba
      1 yersin
      6 yersinia
      3 yerxa
      5 yggdrasil
      1 yijon
      5 yin
      1 ykanaler
      5 ykromosom
      4 ykromosomen
      1 ykromosomer
      1 ykromosomsystem
      1 yled
      2 ylle
      1 yllearbetare
      1 ylletråd
      1 ylletröjor
      2 ylletyger
      2 ymnig
      1 ymnigt
      4 ympning
      2 yngling
      2 ynglingar
      1 ynglingasagan
     61 yngre
      2 yngsta
     59 yoga
      1 yóga
      1 yogafilosofin
      1 yogaläran
      1 yogalärarna
      1 yogametodik
      4 yogan
      2 yogans
      1 yogaövningar
      1 yogarelaterade
      1 yogarörelser
      1 yogaskolan
      1 yogatradition
      1 yogaundervisning
      1 yogautövning
      1 yogendra
      1 yoghurt
      3 yogi
      1 yogini
      1 yōkoso
      1 yolken
     19 york
      2 yorke
      1 yorkshire
      4 you
      1 young
      2 your
      2 youtube
      1 yparametrar
      1 yplattorna
      1 ypperligt
      1 yppigt
      3 yr
      3 yra
      1 yrkade
      1 yrkande
      1 yrkat
     19 yrke
     13 yrken
      1 yrkena
      1 yrkes
      1 yrkesarbetande
      1 yrkesarbetar
      1 yrkesarbete
      1 yrkesbenämningen
      1 yrkesbeteckningen
      2 yrkesbevis
      1 yrkesbeviset
      3 yrkeserfarenhet
      4 yrkesexamen
      1 yrkesexaminan
      1 yrkesförbund
      1 yrkesförbunden
      1 yrkesföreningen
      1 yrkesföreningensveriges
      1 yrkesgrupp
      1 yrkesgruppen
     12 yrkesgrupper
      1 yrkesgrupperna
      1 yrkeshygien
      1 yrkesinriktad
      1 yrkeskår
      2 yrkeskategori
      2 yrkeskategorier
      5 yrkeslegitimation
      1 yrkeslivet
      1 yrkesman
      7 yrkesmässig
      2 yrkesmässiga
      5 yrkesmässigt
      1 yrkesmedicin
      1 yrkesnämnd
      1 yrkesperson
      1 yrkesprofessioner
      1 yrkesprogram
      1 yrkesregister
      1 yrkessjukdom
      2 yrkesskada
      1 yrkesskador
      1 yrkesskyddad
      6 yrkestitel
      5 yrkestiteln
      2 yrkesuppgifter
      5 yrkesutbildning
      1 yrkesutövande
      1 yrkesutövare
      1 yrkesutövningen
      2 yrkesverksam
      2 yrkesverksamhet
      6 yrkesverksamma
      9 yrket
     47 yrsel
      1 yrselförening
      1 yrselpatienter
      1 yrseltillstånd
      1 ysh�ng
      1 yskalan
      1 �ystein
      1 ystenzymer
      1 yt
     46 yta
      1 ytalexi
     25 ytan
      1 ytans
      1 ytarean
      1 ytbehandlade
      1 ytbehandlats
      4 ytbehandling
      1 ytbehandlingsmedel
      3 ytcentrerat
      1 ytdekompression
      1 ytdesinfektion
      2 ytelektroder
      2 ytelektromyografi
      1 ytemg
      1 ytersättning
      1 ytersättningar
      1 ytersättningen
      1 ytersättningsspecialist
      1 ytförstoring
      1 ytkonstruktionen
     13 ytlig
     24 ytliga
      2 ytligare
      8 ytligt
      1 ytmaterial
     16 ytor
      2 ytorna
      3 ytproteiner
      1 ytskikt
      1 ytskrapor
      1 ytslipning
      1 ytspädda
      2 ytspänning
      2 ytstruktur
      1 ytstrukturella
      1 ytstrukturen
      1 ytstrukturerna
      2 ytterdiameter
      1 ytterhölje
      1 ytterjärna
      1 ytterkläder
      1 ytterliga
    162 ytterligare
      1 yttermått
      1 yttermembranet
      1 yttermiljön
      6 ytterörat
      2 ytteröron
      2 ytterplagg
      1 yttersidan
     34 ytterst
     28 yttersta
      1 yttervärlden
     48 yttra
      4 yttrade
      4 yttrande
      1 yttranden
     61 yttrar
    117 yttre
      6 yttringar
      3 ytvatten
      1 ytvattentäkter
      1 yule�walkerekvationerna
      2 yves
      1 yvigare
      1 yvonne
      1 yxa
      1 yxkastning
      4 z
      1 zabern
      1 zacchia
      1 zahra
     13 zaire
      1 zairespecifika
      1 zamiakalla
      1 zamiifolia
      2 zamioculcas
      2 zanamivir
      1 zangwill
      1 zantac
      1 zantedeschia
      1 zanthoxylum
      2 zedrak
     10 zeeland
      1 zeelands
      1 zeiss
      1 zeitgeist
      1 zelmid
      1 zenbuddhismen
      1 zendium
      2 zenker
      1 zetterholm
      1 zetterlund
      2 zeus
      1 zhao
      2 zhongdian
      2 zhou
      1 zhuan
      1 zi
      1 ziehlneelsen
      2 zimbabwe
      3 zimelidin
      1 zinin
     14 zink
      1 zinkånga
      1 zinkblände
      5 zinkbrist
      1 zinkcitrat
      1 zinkfeber
      1 zinkförgiftning
      1 zinkframställningen
      1 zinkfrossa
      1 zinkglukonatpastiller
      2 zinkkarbonat
      1 zinkklorid
      1 zinkkloridkatalysator
      1 zinknivåerna
      3 zinkoxid
      1 zinksulfatlösning
      1 zinksulfid
      2 zinktillskott
      1 zinkvärdena
      1 zinkvitt
      1 zionis
      1 ziprasidon
      2 zkromosom
      1 zkromosomer
      1 zmapp
      3 zo
      1 zodiaken
      9 zolpidem
      1 zolpidems
      2 zon
     19 zona
      1 zonändpunkt
      1 zondek
      1 zone
      2 zonen
      3 zoner
      1 zonlinjer
      1 zonpunkter
      1 zonterapeut
      1 zonterapeuter
      1 zonterapeutiska
      7 zonterapi
      1 zonterapin
      1 zonula
      2 zonulatrådarna
      8 zoo
      1 zoodjur
      1 zooider
      2 zoologen
      2 zoological
      1 zoologiska
      1 zoologiskt
      1 zoology
      1 zoon
     11 zoonos
      1 zoonosa
      4 zoonoser
      6 zoonotisk
      1 zoonotiskt
      1 zoosporer
      1 zootoxin
      2 zoster
      1 zóster
      1 zostervaccination
      3 zostervirus
      1 zovirax
      3 zp
      1 zparametrar
      2 zpglykoproteinerna
      1 zplastik
      1 zscore
     13 zumba
      1 zumbadans
      1 zumbainstruktör
      1 zumban
      1 zumbatomic
      1 zumbaträning
      1 zumbaträningspass
      1 zvärde
      2 zw
      1 zwhonor
      2 zwsystemet
      1 zygosaccharomyces
      4 zygot
      5 zygoten
      1 zygoter
      3 zyklon
      1 zyx
      3 zz
      1 zzbilirubinmolekyl
